

// CBG Orangepath HPR L/S System

// Verilog output file generated at 21/10/2015 18:37:24
// KiwiC (.net/CIL/C# to Verilog/SystemC compiler): Version alpha 56: October-2015 Unix 3.19.8.100
//  /home/djg11/d320/hprls/kiwipro/kiwic/distro/lib/kiwic.exe -verilog-roundtrip=disable -report-each-step -verbose -repack=disable -restructure2=disable sw_test.exe -vnl=disable -sim 100000 -vnl-rootmodname=DUT -kiwic-cil-dump=combined

module DUT(output [31:0] result, output reg signed [63:0] d_monitor, output reg [31:0] phase, input clk, input reset);
  integer TSPru0_12_V_0;
  integer TSPru0_12_V_1;
  integer TSPin0_6_V_0;
  integer TSPen1_8_V_0;
  integer TSPsw1_2_V_0;
  integer TSPsw1_2_V_1;
  integer TSPne2_10_V_0;
  integer TSPne2_10_V_1;
  integer TSPne2_10_V_2;
  integer TSPne2_10_V_3;
  reg signed [63:0] TSPne2_10_V_6;
  integer TSPen0_17_V_0;
  integer TSPte2_13_V_0;
  integer TSPte2_13_V_1;
  integer TSPte2_13_V_2;
  integer TSPcr2_16_V_0;
  integer TSPcr2_16_V_1;
  integer TSPe1_SPILL_256;
  integer TSPe0_SPILL_256;
  reg [9:0] xpc10;
  wire signed [63:0] hprpin256610;
  wire signed [63:0] hprpin258710;
  wire signed [31:0] hprpin529710;
  wire [18:0] hprpin534210;
  wire signed [31:0] hprpin536910;
  wire [18:0] hprpin540610;
 always   @(posedge clk )  begin 
      //Start structure HPR sw_test.exe

      case (xpc10)

      10'd827/*827:US*/: $display("Smith Waterman Simple Test Start. Iterations=%d", 1'd1);

      10'd834/*834:US*/: $display("waypoint %d %d", 2'd2, 0);
      endcase
      if ((32'd1+TSPin0_6_V_0>=7'h4d) && (xpc10==10'd837/*837:US*/)) $display("waypoint %d %d", 2'd3, 0);
          if ((TSPru0_12_V_0>=1'd1) && (xpc10==10'd838/*838:US*/))  begin 
              $display("waypoint %d %d", 4'd12, 0);
              $display("Smith Waterman Simple Test End.");
              $finish(0);
               end 
              if ((TSPru0_12_V_1<7'h4b) && (xpc10==10'd842/*842:US*/))  begin 
              $display("waypoint %d %d", 3'd6, TSPru0_12_V_1);
              $display("waypoint %d %d", 3'd4, 0);
               end 
              if ((TSPne2_10_V_3>=7'h4d) && (xpc10==10'd845/*845:US*/))  begin 
              $display("waypoint %d %d", 4'd8, TSPru0_12_V_1);
              $display("Scored h matrix %d", TSPru0_12_V_1);
               end 
              if ((TSPte2_13_V_0>=2'd2) && (xpc10==10'd846/*846:US*/)) $display("waypoint %d %d", 4'd10, TSPru0_12_V_1);
          if ((TSPcr2_16_V_1>=7'h4d) && (xpc10==10'd847/*847:US*/)) $display("step %d crc is %d", TSPru0_12_V_1, A_UINT[19'h6_3b60+4'd8
          ]);
          
      case (xpc10)

      10'd834/*834:US*/:  begin 
           xpc10 <= 10'd835/*835:xpc10:835*/;
           TSPen1_8_V_0 <= 32'd0;
           TSPin0_6_V_0 <= 32'd0;
           phase <= 32'd2;
           A_SINT[19'h6_353c+4'd8] <= 32'd2;
           end 
          
      10'd837/*837:US*/: if ((32'd1+TSPin0_6_V_0<7'h4d))  begin 
               xpc10 <= 10'd865/*865:xpc10:865*/;
               TSPen1_8_V_0 <= 32'd0;
               TSPin0_6_V_0 <= 32'd1+TSPin0_6_V_0;
               A_SINT[19'h6_3a2c+3'h4*TSPin0_6_V_0] <= TSPe1_SPILL_256;
               end 
               else  begin 
               xpc10 <= 10'd838/*838:xpc10:838*/;
               TSPru0_12_V_0 <= 32'd0;
               phase <= 32'd3;
               TSPin0_6_V_0 <= 32'd1+TSPin0_6_V_0;
               A_SINT[19'h6_3a2c+3'h4*TSPin0_6_V_0] <= TSPe1_SPILL_256;
               end 
              
      10'd838/*838:US*/: if ((TSPru0_12_V_0<1'd1))  xpc10 <= 10'd839/*839:xpc10:839*/;
           else  phase <= 32'd12;

      10'd842/*842:US*/: if ((TSPru0_12_V_1<7'h4b))  begin 
               xpc10 <= 10'd843/*843:xpc10:843*/;
               TSPen0_17_V_0 <= 32'd0;
               TSPne2_10_V_1 <= ((32'd1+TSPru0_12_V_1)%2'd2);
               TSPne2_10_V_0 <= (TSPru0_12_V_1%2'd2);
               phase <= 32'd4;
               end 
               else  begin 
               xpc10 <= 10'd838/*838:xpc10:838*/;
               TSPru0_12_V_0 <= 32'd1+TSPru0_12_V_0;
               end 
              
      10'd845/*845:US*/: if ((TSPne2_10_V_3<7'h4d))  xpc10 <= 10'd850/*850:xpc10:850*/;
           else  begin 
               xpc10 <= 10'd846/*846:xpc10:846*/;
               TSPte2_13_V_0 <= 32'd0;
               phase <= 32'd8+32'd256*TSPru0_12_V_1;
               end 
              
      10'd846/*846:US*/: if ((TSPte2_13_V_0<2'd2))  begin 
               xpc10 <= 10'd848/*848:xpc10:848*/;
               TSPte2_13_V_2 <= 32'd0;
               TSPte2_13_V_1 <= ((TSPru0_12_V_1+TSPte2_13_V_0)%2'd2);
               end 
               else  begin 
               xpc10 <= 10'd847/*847:xpc10:847*/;
               TSPcr2_16_V_1 <= 32'd0;
               TSPcr2_16_V_0 <= ((32'd1+TSPru0_12_V_1)%2'd2);
               phase <= 32'd10+32'd256*TSPru0_12_V_1;
               A_UINT[19'h6_3b60+4'd8] <= -32'd1;
               end 
              
      10'd847/*847:US*/: if ((TSPcr2_16_V_1<7'h4d))  begin 
               TSPcr2_16_V_1 <= 32'd1+TSPcr2_16_V_1;
               A_UINT[19'h6_3b60+4'd8] <= -32'd1&((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c
              +3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))]))? -32'd1&((19'h6_3b60+4'd8==
              19'h6_1a80+3'h4*(8'd255&(hprpin529710>>>5'd16)))? -32'd1&((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255&((-2'd1&A_UINT[19'h6_1a80
              +3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff
              &TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0})>>
              5'd24)))? -32'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff
              &TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24
              ))]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT[32'h6_1a80+3'h4*(8'd255&((-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c
              +4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT
              [19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0})>>5'd24))])^((19'h6_3b60+4'd8
              ==19'h6_1a80+3'h4*(8'd255&(hprpin529710>>>4'd8)))? -32'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT
              [19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80
              +3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT[32'h6_1a80+3'h4*(8'd255&(hprpin529710
              >>>4'd8))])^{-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff
              &TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24
              ))]^{A_UINT[19'h6_3b60+4'd8], 8'd0}, 8'd0}: A_UINT[32'h6_1a80+3'h4*(8'd255&(hprpin529710>>>5'd16))])^((19'h6_3b60+4'd8==
              19'h6_1a80+3'h4*(8'd255&((-2'd1&((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255&((-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS
              [19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1
              ))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0})>>5'd24)))? -32'd1
              &A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0
              )+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT
              [19'h6_3b60+4'd8], 8'd0}: A_UINT[32'h6_1a80+3'h4*(8'd255&((-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8
              *(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80
              +3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0})>>5'd24))])^((19'h6_3b60+4'd8==19'h6_1a80
              +3'h4*(8'd255&(hprpin529710>>>4'd8)))? -32'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c
              +3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255
              &(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT[32'h6_1a80+3'h4*(8'd255&(hprpin529710>>>4'd8
              ))])^{-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0
              )+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT
              [19'h6_3b60+4'd8], 8'd0}, 8'd0})>>5'd24)))? -32'd1&((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255&((-2'd1&A_UINT[19'h6_1a80
              +3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff
              &TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0})>>
              5'd24)))? -32'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff
              &TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24
              ))]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT[32'h6_1a80+3'h4*(8'd255&((-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c
              +4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT
              [19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0})>>5'd24))])^((19'h6_3b60+4'd8
              ==19'h6_1a80+3'h4*(8'd255&(hprpin529710>>>4'd8)))? -32'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT
              [19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80
              +3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT[32'h6_1a80+3'h4*(8'd255&(hprpin529710
              >>>4'd8))])^{-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff
              &TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24
              ))]^{A_UINT[19'h6_3b60+4'd8], 8'd0}, 8'd0}: A_UINT[32'h6_1a80+3'h4*(8'd255&((-2'd1&((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255
              &((-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0
              )+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT
              [19'h6_3b60+4'd8], 8'd0})>>5'd24)))? -32'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4
              ]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&
              (A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT[32'h6_1a80+3'h4*(8'd255&((-2'd1&A_UINT[19'h6_1a80
              +3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff
              &TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0})>>
              5'd24))])^((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255&(hprpin529710>>>4'd8)))? -32'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS
              [19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1
              ))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT[32'h6_1a80
              +3'h4*(8'd255&(hprpin529710>>>4'd8))])^{-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c
              +3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255
              &(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0}, 8'd0})>>5'd24))])^{-2'd1&((19'h6_3b60+4'd8==19'h6_1a80
              +3'h4*(8'd255&((-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff
              &TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24
              ))]^{A_UINT[19'h6_3b60+4'd8], 8'd0})>>5'd24)))? -32'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c
              +3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255
              &(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT[32'h6_1a80+3'h4*(8'd255&((-2'd1&A_UINT[19'h6_1a80
              +3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff
              &TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0})>>
              5'd24))])^((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255&(hprpin529710>>>4'd8)))? -32'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS
              [19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1
              ))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT[32'h6_1a80
              +3'h4*(8'd255&(hprpin529710>>>4'd8))])^{-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c
              +3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255
              &(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0}, 8'd0}, 8'd0}: A_UINT[32'h6_1a80+3'h4*(8'd255&A_64_SS
              [19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1
              ))])])^((hprpin534210==19'h6_3b60+4'd8)? -32'd1&((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255&(hprpin529710>>>5'd16)))? -32'd1
              &((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255&((-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c
              +3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255
              &(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0})>>5'd24)))? -32'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS
              [19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1
              ))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT[32'h6_1a80
              +3'h4*(8'd255&((-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff
              &TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24
              ))]^{A_UINT[19'h6_3b60+4'd8], 8'd0})>>5'd24))])^((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255&(hprpin529710>>>4'd8)))? -32'd1
              &A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0
              )+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT
              [19'h6_3b60+4'd8], 8'd0}: A_UINT[32'h6_1a80+3'h4*(8'd255&(hprpin529710>>>4'd8))])^{-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255
              &A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1
              ))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0}, 8'd0}: A_UINT[32'h6_1a80
              +3'h4*(8'd255&(hprpin529710>>>5'd16))])^((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255&((-2'd1&((19'h6_3b60+4'd8==19'h6_1a80
              +3'h4*(8'd255&((-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff
              &TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24
              ))]^{A_UINT[19'h6_3b60+4'd8], 8'd0})>>5'd24)))? -32'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c
              +3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255
              &(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT[32'h6_1a80+3'h4*(8'd255&((-2'd1&A_UINT[19'h6_1a80
              +3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff
              &TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0})>>
              5'd24))])^((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255&(hprpin529710>>>4'd8)))? -32'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS
              [19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1
              ))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT[32'h6_1a80
              +3'h4*(8'd255&(hprpin529710>>>4'd8))])^{-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c
              +3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255
              &(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0}, 8'd0})>>5'd24)))? -32'd1&((19'h6_3b60+4'd8==19'h6_1a80
              +3'h4*(8'd255&((-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff
              &TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24
              ))]^{A_UINT[19'h6_3b60+4'd8], 8'd0})>>5'd24)))? -32'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c
              +3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255
              &(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT[32'h6_1a80+3'h4*(8'd255&((-2'd1&A_UINT[19'h6_1a80
              +3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff
              &TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0})>>
              5'd24))])^((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255&(hprpin529710>>>4'd8)))? -32'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS
              [19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1
              ))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT[32'h6_1a80
              +3'h4*(8'd255&(hprpin529710>>>4'd8))])^{-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c
              +3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255
              &(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0}, 8'd0}: A_UINT[32'h6_1a80+3'h4*(8'd255&((-2'd1&((19'h6_3b60
              +4'd8==19'h6_1a80+3'h4*(8'd255&((-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*
              (64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT
              [19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0})>>5'd24)))? -32'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c
              +4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT
              [19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT[32'h6_1a80+3'h4*(8'd255
              &((-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0
              )+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT
              [19'h6_3b60+4'd8], 8'd0})>>5'd24))])^((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255&(hprpin529710>>>4'd8)))? -32'd1&A_UINT[19'h6_1a80
              +3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff
              &TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT
              [32'h6_1a80+3'h4*(8'd255&(hprpin529710>>>4'd8))])^{-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT
              [19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80
              +3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0}, 8'd0})>>5'd24))])^{-2'd1&((19'h6_3b60
              +4'd8==19'h6_1a80+3'h4*(8'd255&((-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*
              (64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT
              [19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0})>>5'd24)))? -32'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c
              +4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT
              [19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT[32'h6_1a80+3'h4*(8'd255
              &((-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0
              )+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT
              [19'h6_3b60+4'd8], 8'd0})>>5'd24))])^((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255&(hprpin529710>>>4'd8)))? -32'd1&A_UINT[19'h6_1a80
              +3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff
              &TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT
              [32'h6_1a80+3'h4*(8'd255&(hprpin529710>>>4'd8))])^{-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT
              [19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80
              +3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0}, 8'd0}, 8'd0}: A_UINT[hprpin534210])^{-32'd1
              &((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255&(hprpin529710>>>5'd16)))? -32'd1&((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255
              &((-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0
              )+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT
              [19'h6_3b60+4'd8], 8'd0})>>5'd24)))? -32'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4
              ]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&
              (A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT[32'h6_1a80+3'h4*(8'd255&((-2'd1&A_UINT[19'h6_1a80
              +3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff
              &TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0})>>
              5'd24))])^((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255&(hprpin529710>>>4'd8)))? -32'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS
              [19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1
              ))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT[32'h6_1a80
              +3'h4*(8'd255&(hprpin529710>>>4'd8))])^{-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c
              +3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255
              &(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0}, 8'd0}: A_UINT[32'h6_1a80+3'h4*(8'd255&(hprpin529710
              >>>5'd16))])^((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255&((-2'd1&((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255&((-2'd1&A_UINT
              [19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff
              &TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0})>>
              5'd24)))? -32'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff
              &TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24
              ))]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT[32'h6_1a80+3'h4*(8'd255&((-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c
              +4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT
              [19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0})>>5'd24))])^((19'h6_3b60+4'd8
              ==19'h6_1a80+3'h4*(8'd255&(hprpin529710>>>4'd8)))? -32'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT
              [19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80
              +3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT[32'h6_1a80+3'h4*(8'd255&(hprpin529710
              >>>4'd8))])^{-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff
              &TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24
              ))]^{A_UINT[19'h6_3b60+4'd8], 8'd0}, 8'd0})>>5'd24)))? -32'd1&((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255&((-2'd1&A_UINT
              [19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff
              &TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0})>>
              5'd24)))? -32'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff
              &TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24
              ))]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT[32'h6_1a80+3'h4*(8'd255&((-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c
              +4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT
              [19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0})>>5'd24))])^((19'h6_3b60+4'd8
              ==19'h6_1a80+3'h4*(8'd255&(hprpin529710>>>4'd8)))? -32'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT
              [19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80
              +3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT[32'h6_1a80+3'h4*(8'd255&(hprpin529710
              >>>4'd8))])^{-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff
              &TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24
              ))]^{A_UINT[19'h6_3b60+4'd8], 8'd0}, 8'd0}: A_UINT[32'h6_1a80+3'h4*(8'd255&((-2'd1&((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255
              &((-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0
              )+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT
              [19'h6_3b60+4'd8], 8'd0})>>5'd24)))? -32'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4
              ]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&
              (A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT[32'h6_1a80+3'h4*(8'd255&((-2'd1&A_UINT[19'h6_1a80
              +3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff
              &TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0})>>
              5'd24))])^((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255&(hprpin529710>>>4'd8)))? -32'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS
              [19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1
              ))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT[32'h6_1a80
              +3'h4*(8'd255&(hprpin529710>>>4'd8))])^{-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c
              +3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255
              &(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0}, 8'd0})>>5'd24))])^{-2'd1&((19'h6_3b60+4'd8==19'h6_1a80
              +3'h4*(8'd255&((-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff
              &TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24
              ))]^{A_UINT[19'h6_3b60+4'd8], 8'd0})>>5'd24)))? -32'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c
              +3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255
              &(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT[32'h6_1a80+3'h4*(8'd255&((-2'd1&A_UINT[19'h6_1a80
              +3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff
              &TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0})>>
              5'd24))])^((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255&(hprpin529710>>>4'd8)))? -32'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS
              [19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1
              ))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT[32'h6_1a80
              +3'h4*(8'd255&(hprpin529710>>>4'd8))])^{-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c
              +3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255
              &(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0}, 8'd0}, 8'd0}, 8'd0};

               end 
               else  begin 
               xpc10 <= 10'd842/*842:xpc10:842*/;
               TSPru0_12_V_1 <= 32'd1+TSPru0_12_V_1;
               d_monitor <= 64'h_ffff_ffff_ffff_ffff&A_UINT[19'h6_3b60+4'd8];
               end 
              
      10'd849/*849:US*/:  begin 
          $write("%d %d : %d   ", TSPte2_13_V_1, TSPte2_13_V_2, A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff
          &TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))]);
          $display("");
           xpc10 <= 10'd848/*848:xpc10:848*/;
           TSPte2_13_V_2 <= 32'd1+TSPte2_13_V_2;
           A_UINT[19'h6_3b60+4'd8] <= -32'd1&((hprpin540610==19'h6_3b60+4'd8)? -32'd1&((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255&((-2'd1
          &((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255&((-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT
          [19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff
          &TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0})>>5'd24)))? -2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8
          ]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1
          )+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT[19'h6_1a80+3'h4*(8'd255&((-2'd1&A_UINT
          [19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c
          +3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0
          })>>5'd24))])^((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255&(hprpin536910>>>4'd8)))? -2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT
          [19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff
          &TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT[19'h6_1a80+3'h4*(8'd255
          &(hprpin536910>>>4'd8))])^{-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255
          &A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2
          ))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0}, 8'd0})>>5'd24)))? -32'd1&((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255&((-2'd1&A_UINT[19'h6_1a80
          +3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+
          3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0})>>
          5'd24)))? -2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c
          +4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT
          [19'h6_3b60+4'd8], 8'd0}: A_UINT[19'h6_1a80+3'h4*(8'd255&((-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24
          ))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1
          )+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0})>>5'd24))])^((19'h6_3b60+4'd8==19'h6_1a80+3'h4
          *(8'd255&(hprpin536910>>>4'd8)))? -2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80
          +3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff
          &TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT[19'h6_1a80+3'h4*(8'd255&(hprpin536910>>>4'd8))])^{-2'd1&A_UINT[19'h6_1a80
          +3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+
          3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0}, 8'd0
          }: A_UINT[32'h6_1a80+3'h4*(8'd255&((-2'd1&((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255&((-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255
          &(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff
          &TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0})>>5'd24)))? -2'd1&A_UINT[19'h6_1a80
          +3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+
          3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT
          [19'h6_1a80+3'h4*(8'd255&((-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255
          &A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2
          ))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0})>>5'd24))])^((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255&(hprpin536910>>>4'd8)))? -2'd1
          &A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT
          [19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+
          4'd8], 8'd0}: A_UINT[19'h6_1a80+3'h4*(8'd255&(hprpin536910>>>4'd8))])^{-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60
          +4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&
          TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0}, 8'd0})>>5'd24))])^((19'h6_3b60
          +4'd8==19'h6_1a80+3'h4*(8'd255&(hprpin536910>>>5'd16)))? -32'd1&((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255&((-2'd1&A_UINT[19'h6_1a80
          +3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+
          3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0})>>
          5'd24)))? -2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c
          +4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT
          [19'h6_3b60+4'd8], 8'd0}: A_UINT[19'h6_1a80+3'h4*(8'd255&((-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24
          ))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1
          )+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0})>>5'd24))])^((19'h6_3b60+4'd8==19'h6_1a80+3'h4
          *(8'd255&(hprpin536910>>>4'd8)))? -2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80
          +3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff
          &TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT[19'h6_1a80+3'h4*(8'd255&(hprpin536910>>>4'd8))])^{-2'd1&A_UINT[19'h6_1a80
          +3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+
          3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0}, 8'd0
          }: A_UINT[32'h6_1a80+3'h4*(8'd255&(hprpin536910>>>5'd16))])^{-2'd1&((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255&((-2'd1&A_UINT
          [19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c
          +3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0
          })>>5'd24)))? -2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS
          [19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))]
          )]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT[19'h6_1a80+3'h4*(8'd255&((-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60
          +4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&
          TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0})>>5'd24))])^((19'h6_3b60+4'd8==
          19'h6_1a80+3'h4*(8'd255&(hprpin536910>>>4'd8)))? -2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT
          [19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff
          &TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT[19'h6_1a80+3'h4*(8'd255&(hprpin536910>>>4'd8))])^{-2'd1&A_UINT[19'h6_1a80
          +3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+
          3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0}, 8'd0
          }, 8'd0}: A_UINT[hprpin540610])^((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]
          *(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))]))? -32'd1&((19'h6_3b60+4'd8==19'h6_1a80
          +3'h4*(8'd255&((-2'd1&((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255&((-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+
          4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1
          )+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0})>>5'd24)))? -2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255
          &(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff
          &TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT[19'h6_1a80+3'h4*(8'd255
          &((-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c
          +4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT
          [19'h6_3b60+4'd8], 8'd0})>>5'd24))])^((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255&(hprpin536910>>>4'd8)))? -2'd1&A_UINT[19'h6_1a80
          +3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+
          3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT
          [19'h6_1a80+3'h4*(8'd255&(hprpin536910>>>4'd8))])^{-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^
          A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff
          &TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0}, 8'd0})>>5'd24)))? -32'd1&((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255&((-2'd1
          &A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT
          [19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+
          4'd8], 8'd0})>>5'd24)))? -2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255
          &A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2
          ))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT[19'h6_1a80+3'h4*(8'd255&((-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60
          +4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&
          TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0})>>5'd24))])^((19'h6_3b60+4'd8==
          19'h6_1a80+3'h4*(8'd255&(hprpin536910>>>4'd8)))? -2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT
          [19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff
          &TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT[19'h6_1a80+3'h4*(8'd255&(hprpin536910>>>4'd8))])^{-2'd1&A_UINT[19'h6_1a80
          +3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+
          3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0}, 8'd0
          }: A_UINT[32'h6_1a80+3'h4*(8'd255&((-2'd1&((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255&((-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255
          &(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff
          &TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0})>>5'd24)))? -2'd1&A_UINT[19'h6_1a80
          +3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+
          3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT
          [19'h6_1a80+3'h4*(8'd255&((-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255
          &A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2
          ))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0})>>5'd24))])^((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255&(hprpin536910>>>4'd8)))? -2'd1
          &A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT
          [19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+
          4'd8], 8'd0}: A_UINT[19'h6_1a80+3'h4*(8'd255&(hprpin536910>>>4'd8))])^{-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60
          +4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&
          TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0}, 8'd0})>>5'd24))])^((19'h6_3b60
          +4'd8==19'h6_1a80+3'h4*(8'd255&(hprpin536910>>>5'd16)))? -32'd1&((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255&((-2'd1&A_UINT[19'h6_1a80
          +3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+
          3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0})>>
          5'd24)))? -2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c
          +4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT
          [19'h6_3b60+4'd8], 8'd0}: A_UINT[19'h6_1a80+3'h4*(8'd255&((-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24
          ))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1
          )+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0})>>5'd24))])^((19'h6_3b60+4'd8==19'h6_1a80+3'h4
          *(8'd255&(hprpin536910>>>4'd8)))? -2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80
          +3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff
          &TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT[19'h6_1a80+3'h4*(8'd255&(hprpin536910>>>4'd8))])^{-2'd1&A_UINT[19'h6_1a80
          +3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+
          3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0}, 8'd0
          }: A_UINT[32'h6_1a80+3'h4*(8'd255&(hprpin536910>>>5'd16))])^{-2'd1&((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255&((-2'd1&A_UINT
          [19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c
          +3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0
          })>>5'd24)))? -2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS
          [19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))]
          )]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT[19'h6_1a80+3'h4*(8'd255&((-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60
          +4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&
          TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0})>>5'd24))])^((19'h6_3b60+4'd8==
          19'h6_1a80+3'h4*(8'd255&(hprpin536910>>>4'd8)))? -2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT
          [19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff
          &TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT[19'h6_1a80+3'h4*(8'd255&(hprpin536910>>>4'd8))])^{-2'd1&A_UINT[19'h6_1a80
          +3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+
          3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0}, 8'd0
          }, 8'd0}: A_UINT[32'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1
          )+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])])^{-32'd1&((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255&((-2'd1&((19'h6_3b60+4'd8
          ==19'h6_1a80+3'h4*(8'd255&((-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*
          (8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff
          &TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0})>>5'd24)))? -2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8
          ]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1
          )+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT[19'h6_1a80+3'h4*(8'd255&((-2'd1&A_UINT
          [19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c
          +3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0
          })>>5'd24))])^((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255&(hprpin536910>>>4'd8)))? -2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT
          [19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff
          &TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT[19'h6_1a80+3'h4*(8'd255
          &(hprpin536910>>>4'd8))])^{-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255
          &A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2
          ))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0}, 8'd0})>>5'd24)))? -32'd1&((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255&((-2'd1&A_UINT[19'h6_1a80
          +3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+
          3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0})>>
          5'd24)))? -2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c
          +4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT
          [19'h6_3b60+4'd8], 8'd0}: A_UINT[19'h6_1a80+3'h4*(8'd255&((-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24
          ))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1
          )+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0})>>5'd24))])^((19'h6_3b60+4'd8==19'h6_1a80+3'h4
          *(8'd255&(hprpin536910>>>4'd8)))? -2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80
          +3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff
          &TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT[19'h6_1a80+3'h4*(8'd255&(hprpin536910>>>4'd8))])^{-2'd1&A_UINT[19'h6_1a80
          +3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+
          3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0}, 8'd0
          }: A_UINT[32'h6_1a80+3'h4*(8'd255&((-2'd1&((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255&((-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255
          &(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff
          &TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0})>>5'd24)))? -2'd1&A_UINT[19'h6_1a80
          +3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+
          3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT
          [19'h6_1a80+3'h4*(8'd255&((-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255
          &A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2
          ))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0})>>5'd24))])^((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255&(hprpin536910>>>4'd8)))? -2'd1
          &A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT
          [19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+
          4'd8], 8'd0}: A_UINT[19'h6_1a80+3'h4*(8'd255&(hprpin536910>>>4'd8))])^{-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60
          +4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&
          TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0}, 8'd0})>>5'd24))])^((19'h6_3b60
          +4'd8==19'h6_1a80+3'h4*(8'd255&(hprpin536910>>>5'd16)))? -32'd1&((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255&((-2'd1&A_UINT[19'h6_1a80
          +3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+
          3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0})>>
          5'd24)))? -2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c
          +4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT
          [19'h6_3b60+4'd8], 8'd0}: A_UINT[19'h6_1a80+3'h4*(8'd255&((-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24
          ))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1
          )+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0})>>5'd24))])^((19'h6_3b60+4'd8==19'h6_1a80+3'h4
          *(8'd255&(hprpin536910>>>4'd8)))? -2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80
          +3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff
          &TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT[19'h6_1a80+3'h4*(8'd255&(hprpin536910>>>4'd8))])^{-2'd1&A_UINT[19'h6_1a80
          +3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+
          3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0}, 8'd0
          }: A_UINT[32'h6_1a80+3'h4*(8'd255&(hprpin536910>>>5'd16))])^{-2'd1&((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255&((-2'd1&A_UINT
          [19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c
          +3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0
          })>>5'd24)))? -2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS
          [19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))]
          )]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT[19'h6_1a80+3'h4*(8'd255&((-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60
          +4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&
          TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0})>>5'd24))])^((19'h6_3b60+4'd8==
          19'h6_1a80+3'h4*(8'd255&(hprpin536910>>>4'd8)))? -2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT
          [19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff
          &TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT[19'h6_1a80+3'h4*(8'd255&(hprpin536910>>>4'd8))])^{-2'd1&A_UINT[19'h6_1a80
          +3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+
          3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0}, 8'd0
          }, 8'd0}, 8'd0};

           end 
          endcase
      if ((A_16_SS[19'h6_1f42+2'h2*TSPru0_12_V_1]==A_16_SS[19'h6_1e80+2'h2*TSPen0_17_V_0]))  begin if ((xpc10==10'd856/*856:US*/))  begin 
                   xpc10 <= 10'd844/*844:xpc10:844*/;
                   TSPe0_SPILL_256 <= TSPen0_17_V_0;
                   end 
                   end 
           else if ((xpc10==10'd856/*856:US*/))  begin 
                   xpc10 <= 10'd843/*843:xpc10:843*/;
                   TSPen0_17_V_0 <= 32'd1+TSPen0_17_V_0;
                   end 
                  
      case (xpc10)

      10'd850/*850:US*/: if ((-64'd2+A_64_SS[64'h6_267c+64'h8*(A_SINT[19'h6_266c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPne2_10_V_0)+(64'h_ffff_ffff_ffff_ffff
      &1'd1+TSPne2_10_V_3))]<A_64_SS[19'h6_354c+4'h8*(A_SINT[19'h6_353c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPne2_10_V_0)+(64'h_ffff_ffff_ffff_ffff
      &1'd1+TSPne2_10_V_3))]))  begin 
               xpc10 <= 10'd851/*851:xpc10:851*/;
               A_64_SS[19'h6_267c+4'h8*(A_SINT[19'h6_266c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPne2_10_V_1)+(64'h_ffff_ffff_ffff_ffff&1'd1
              +TSPne2_10_V_3))] <= hprpin256610;

               end 
               else  begin 
               xpc10 <= 10'd851/*851:xpc10:851*/;
               A_64_SS[19'h6_267c+4'h8*(A_SINT[19'h6_266c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPne2_10_V_1)+(64'h_ffff_ffff_ffff_ffff&1'd1
              +TSPne2_10_V_3))] <= -64'd2+A_64_SS[64'h6_267c+64'h8*(A_SINT[19'h6_266c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPne2_10_V_0)+
              (64'h_ffff_ffff_ffff_ffff&1'd1+TSPne2_10_V_3))];

               end 
              
      10'd851/*851:US*/: if ((-3'd2+A_64_SS[19'h6_2b6c+4'h8*(A_SINT[19'h6_2b5c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPne2_10_V_1)+(64'h_ffff_ffff_ffff_ffff
      &TSPne2_10_V_3))]<A_64_SS[64'h6_354c+64'h8*(A_SINT[19'h6_353c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPne2_10_V_1)+(64'h_ffff_ffff_ffff_ffff
      &TSPne2_10_V_3))]))  begin 
               xpc10 <= 10'd852/*852:xpc10:852*/;
               A_64_SS[19'h6_2b6c+4'h8*(A_SINT[19'h6_2b5c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPne2_10_V_1)+(64'h_ffff_ffff_ffff_ffff&1'd1
              +TSPne2_10_V_3))] <= A_64_SS[64'h6_354c+64'h8*(A_SINT[19'h6_353c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPne2_10_V_1)+(64'h_ffff_ffff_ffff_ffff
              &TSPne2_10_V_3))];

               end 
               else  begin 
               xpc10 <= 10'd852/*852:xpc10:852*/;
               A_64_SS[19'h6_267c+4'h8*(A_SINT[19'h6_266c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPne2_10_V_1)+(64'h_ffff_ffff_ffff_ffff&1'd1
              +TSPne2_10_V_3))] <= hprpin258710;

               end 
              
      10'd852/*852:US*/: if ((A_64_SS[64'h6_2b6c+64'h8*(A_SINT[19'h6_2b5c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPne2_10_V_0)+(64'h_ffff_ffff_ffff_ffff
      &TSPne2_10_V_3))]<A_64_SS[64'h6_267c+64'h8*(A_SINT[19'h6_266c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPne2_10_V_0)+(64'h_ffff_ffff_ffff_ffff
      &TSPne2_10_V_3))]))  begin 
               xpc10 <= 10'd853/*853:xpc10:853*/;
               TSPne2_10_V_6 <= A_64_SS[64'h6_267c+64'h8*(A_SINT[19'h6_266c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPne2_10_V_0)+(64'h_ffff_ffff_ffff_ffff
              &TSPne2_10_V_3))];

               end 
               else  begin 
               xpc10 <= 10'd853/*853:xpc10:853*/;
               TSPne2_10_V_6 <= A_64_SS[64'h6_2b6c+64'h8*(A_SINT[19'h6_2b5c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPne2_10_V_0)+(64'h_ffff_ffff_ffff_ffff
              &TSPne2_10_V_3))];

               end 
              
      10'd854/*854:US*/: if ((A_SINT[64'h6_1fe8+64'h4*(A_SINT[64'h6_1fd8+64'd4]*(64'h_ffff_ffff_ffff_ffff&A_SINT[64'h6_3a2c+64'h4*TSPne2_10_V_3
      ])+(64'h_ffff_ffff_ffff_ffff&TSPne2_10_V_2))]+TSPne2_10_V_6<0))  begin 
               xpc10 <= 10'd855/*855:xpc10:855*/;
               A_64_SS[64'h6_305c+64'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPne2_10_V_1)+(64'h_ffff_ffff_ffff_ffff&1'd1
              +TSPne2_10_V_3))] <= 64'd0;

               end 
               else  begin 
               xpc10 <= 10'd855/*855:xpc10:855*/;
               A_64_SS[64'h6_305c+64'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPne2_10_V_1)+(64'h_ffff_ffff_ffff_ffff&1'd1
              +TSPne2_10_V_3))] <= A_SINT[64'h6_1fe8+64'h4*(A_SINT[64'h6_1fd8+64'd4]*(64'h_ffff_ffff_ffff_ffff&A_SINT[64'h6_3a2c+64'h4
              *TSPne2_10_V_3])+(64'h_ffff_ffff_ffff_ffff&TSPne2_10_V_2))]+TSPne2_10_V_6;

               end 
              endcase
      if ((A_16_SS[19'h6_1ea8+2'h2*TSPin0_6_V_0]==A_16_SS[19'h6_1e80+2'h2*TSPen1_8_V_0]))  begin if ((xpc10==10'd836/*836:US*/))  begin 
                   xpc10 <= 10'd837/*837:xpc10:837*/;
                   TSPe1_SPILL_256 <= TSPen1_8_V_0;
                   end 
                   end 
           else if ((xpc10==10'd836/*836:US*/))  begin 
                   xpc10 <= 10'd865/*865:xpc10:865*/;
                   TSPen1_8_V_0 <= 32'd1+TSPen1_8_V_0;
                   end 
                  
      case (xpc10)

      0/*0:US*/:  begin 
           xpc10 <= 1'd1/*1:xpc10:1*/;
           A_16_SS[19'h6_1e80+0] <= 16'd97;
           end 
          
      1'd1/*1:US*/:  begin 
           xpc10 <= 2'd2/*2:xpc10:2*/;
           A_16_SS[19'h6_1e80+2'h2] <= 16'd99;
           end 
          
      2'd2/*2:US*/:  begin 
           xpc10 <= 2'd3/*3:xpc10:3*/;
           A_16_SS[19'h6_1e80+3'h4] <= 16'd100;
           end 
          
      2'd3/*3:US*/:  begin 
           xpc10 <= 3'd4/*4:xpc10:4*/;
           A_16_SS[19'h6_1e80+3'h6] <= 16'd101;
           end 
          
      3'd4/*4:US*/:  begin 
           xpc10 <= 3'd5/*5:xpc10:5*/;
           A_16_SS[19'h6_1e80+4'h8] <= 16'd102;
           end 
          
      3'd5/*5:US*/:  begin 
           xpc10 <= 3'd6/*6:xpc10:6*/;
           A_16_SS[19'h6_1e80+4'ha] <= 16'd103;
           end 
          
      3'd6/*6:US*/:  begin 
           xpc10 <= 3'd7/*7:xpc10:7*/;
           A_16_SS[19'h6_1e80+4'hc] <= 16'd104;
           end 
          
      3'd7/*7:US*/:  begin 
           xpc10 <= 4'd8/*8:xpc10:8*/;
           A_16_SS[19'h6_1e80+4'he] <= 16'd105;
           end 
          
      4'd8/*8:US*/:  begin 
           xpc10 <= 4'd9/*9:xpc10:9*/;
           A_16_SS[19'h6_1e80+5'h10] <= 16'd107;
           end 
          
      4'd9/*9:US*/:  begin 
           xpc10 <= 4'd10/*10:xpc10:10*/;
           A_16_SS[19'h6_1e80+5'h12] <= 16'd108;
           end 
          
      4'd10/*10:US*/:  begin 
           xpc10 <= 4'd11/*11:xpc10:11*/;
           A_16_SS[19'h6_1e80+5'h14] <= 16'd109;
           end 
          
      4'd11/*11:US*/:  begin 
           xpc10 <= 4'd12/*12:xpc10:12*/;
           A_16_SS[19'h6_1e80+5'h16] <= 16'd110;
           end 
          
      4'd12/*12:US*/:  begin 
           xpc10 <= 4'd13/*13:xpc10:13*/;
           A_16_SS[19'h6_1e80+5'h18] <= 16'd112;
           end 
          
      4'd13/*13:US*/:  begin 
           xpc10 <= 4'd14/*14:xpc10:14*/;
           A_16_SS[19'h6_1e80+5'h1a] <= 16'd113;
           end 
          
      4'd14/*14:US*/:  begin 
           xpc10 <= 4'd15/*15:xpc10:15*/;
           A_16_SS[19'h6_1e80+5'h1c] <= 16'd114;
           end 
          
      4'd15/*15:US*/:  begin 
           xpc10 <= 5'd16/*16:xpc10:16*/;
           A_16_SS[19'h6_1e80+5'h1e] <= 16'd115;
           end 
          
      5'd16/*16:US*/:  begin 
           xpc10 <= 5'd17/*17:xpc10:17*/;
           A_16_SS[19'h6_1e80+6'h20] <= 16'd116;
           end 
          
      5'd17/*17:US*/:  begin 
           xpc10 <= 5'd18/*18:xpc10:18*/;
           A_16_SS[19'h6_1e80+6'h22] <= 16'd118;
           end 
          
      5'd18/*18:US*/:  begin 
           xpc10 <= 5'd19/*19:xpc10:19*/;
           A_16_SS[19'h6_1e80+6'h24] <= 16'd119;
           end 
          
      5'd19/*19:US*/:  begin 
           xpc10 <= 5'd20/*20:xpc10:20*/;
           A_16_SS[19'h6_1e80+6'h26] <= 16'd121;
           end 
          
      5'd20/*20:US*/:  begin 
           xpc10 <= 5'd21/*21:xpc10:21*/;
           A_16_SS[19'h6_1ea8+0] <= 16'd100;
           end 
          
      5'd21/*21:US*/:  begin 
           xpc10 <= 5'd22/*22:xpc10:22*/;
           A_16_SS[19'h6_1ea8+2'h2] <= 16'd107;
           end 
          
      5'd22/*22:US*/:  begin 
           xpc10 <= 5'd23/*23:xpc10:23*/;
           A_16_SS[19'h6_1ea8+3'h4] <= 16'd104;
           end 
          
      5'd23/*23:US*/:  begin 
           xpc10 <= 5'd24/*24:xpc10:24*/;
           A_16_SS[19'h6_1ea8+3'h6] <= 16'd107;
           end 
          
      5'd24/*24:US*/:  begin 
           xpc10 <= 5'd25/*25:xpc10:25*/;
           A_16_SS[19'h6_1ea8+4'h8] <= 16'd108;
           end 
          
      5'd25/*25:US*/:  begin 
           xpc10 <= 5'd26/*26:xpc10:26*/;
           A_16_SS[19'h6_1ea8+4'ha] <= 16'd105;
           end 
          
      5'd26/*26:US*/:  begin 
           xpc10 <= 5'd27/*27:xpc10:27*/;
           A_16_SS[19'h6_1ea8+4'hc] <= 16'd116;
           end 
          
      5'd27/*27:US*/:  begin 
           xpc10 <= 5'd28/*28:xpc10:28*/;
           A_16_SS[19'h6_1ea8+4'he] <= 16'd107;
           end 
          
      5'd28/*28:US*/:  begin 
           xpc10 <= 5'd29/*29:xpc10:29*/;
           A_16_SS[19'h6_1ea8+5'h10] <= 16'd116;
           end 
          
      5'd29/*29:US*/:  begin 
           xpc10 <= 5'd30/*30:xpc10:30*/;
           A_16_SS[19'h6_1ea8+5'h12] <= 16'd101;
           end 
          
      5'd30/*30:US*/:  begin 
           xpc10 <= 5'd31/*31:xpc10:31*/;
           A_16_SS[19'h6_1ea8+5'h14] <= 16'd97;
           end 
          
      5'd31/*31:US*/:  begin 
           xpc10 <= 6'd32/*32:xpc10:32*/;
           A_16_SS[19'h6_1ea8+5'h16] <= 16'd107;
           end 
          
      6'd32/*32:US*/:  begin 
           xpc10 <= 6'd33/*33:xpc10:33*/;
           A_16_SS[19'h6_1ea8+5'h18] <= 16'd113;
           end 
          
      6'd33/*33:US*/:  begin 
           xpc10 <= 6'd34/*34:xpc10:34*/;
           A_16_SS[19'h6_1ea8+5'h1a] <= 16'd101;
           end 
          
      6'd34/*34:US*/:  begin 
           xpc10 <= 6'd35/*35:xpc10:35*/;
           A_16_SS[19'h6_1ea8+5'h1c] <= 16'd121;
           end 
          
      6'd35/*35:US*/:  begin 
           xpc10 <= 6'd36/*36:xpc10:36*/;
           A_16_SS[19'h6_1ea8+5'h1e] <= 16'd108;
           end 
          
      6'd36/*36:US*/:  begin 
           xpc10 <= 6'd37/*37:xpc10:37*/;
           A_16_SS[19'h6_1ea8+6'h20] <= 16'd108;
           end 
          
      6'd37/*37:US*/:  begin 
           xpc10 <= 6'd38/*38:xpc10:38*/;
           A_16_SS[19'h6_1ea8+6'h22] <= 16'd107;
           end 
          
      6'd38/*38:US*/:  begin 
           xpc10 <= 6'd39/*39:xpc10:39*/;
           A_16_SS[19'h6_1ea8+6'h24] <= 16'd100;
           end 
          
      6'd39/*39:US*/:  begin 
           xpc10 <= 6'd40/*40:xpc10:40*/;
           A_16_SS[19'h6_1ea8+6'h26] <= 16'd99;
           end 
          
      6'd40/*40:US*/:  begin 
           xpc10 <= 6'd41/*41:xpc10:41*/;
           A_16_SS[19'h6_1ea8+6'h28] <= 16'd100;
           end 
          
      6'd41/*41:US*/:  begin 
           xpc10 <= 6'd42/*42:xpc10:42*/;
           A_16_SS[19'h6_1ea8+6'h2a] <= 16'd108;
           end 
          
      6'd42/*42:US*/:  begin 
           xpc10 <= 6'd43/*43:xpc10:43*/;
           A_16_SS[19'h6_1ea8+6'h2c] <= 16'd101;
           end 
          
      6'd43/*43:US*/:  begin 
           xpc10 <= 6'd44/*44:xpc10:44*/;
           A_16_SS[19'h6_1ea8+6'h2e] <= 16'd107;
           end 
          
      6'd44/*44:US*/:  begin 
           xpc10 <= 6'd45/*45:xpc10:45*/;
           A_16_SS[19'h6_1ea8+6'h30] <= 16'd114;
           end 
          
      6'd45/*45:US*/:  begin 
           xpc10 <= 6'd46/*46:xpc10:46*/;
           A_16_SS[19'h6_1ea8+6'h32] <= 16'd101;
           end 
          
      6'd46/*46:US*/:  begin 
           xpc10 <= 6'd47/*47:xpc10:47*/;
           A_16_SS[19'h6_1ea8+6'h34] <= 16'd112;
           end 
          
      6'd47/*47:US*/:  begin 
           xpc10 <= 6'd48/*48:xpc10:48*/;
           A_16_SS[19'h6_1ea8+6'h36] <= 16'd112;
           end 
          
      6'd48/*48:US*/:  begin 
           xpc10 <= 6'd49/*49:xpc10:49*/;
           A_16_SS[19'h6_1ea8+6'h38] <= 16'd108;
           end 
          
      6'd49/*49:US*/:  begin 
           xpc10 <= 6'd50/*50:xpc10:50*/;
           A_16_SS[19'h6_1ea8+6'h3a] <= 16'd107;
           end 
          
      6'd50/*50:US*/:  begin 
           xpc10 <= 6'd51/*51:xpc10:51*/;
           A_16_SS[19'h6_1ea8+6'h3c] <= 16'd102;
           end 
          
      6'd51/*51:US*/:  begin 
           xpc10 <= 6'd52/*52:xpc10:52*/;
           A_16_SS[19'h6_1ea8+6'h3e] <= 16'd105;
           end 
          
      6'd52/*52:US*/:  begin 
           xpc10 <= 6'd53/*53:xpc10:53*/;
           A_16_SS[19'h6_1ea8+7'h40] <= 16'd118;
           end 
          
      6'd53/*53:US*/:  begin 
           xpc10 <= 6'd54/*54:xpc10:54*/;
           A_16_SS[19'h6_1ea8+7'h42] <= 16'd107;
           end 
          
      6'd54/*54:US*/:  begin 
           xpc10 <= 6'd55/*55:xpc10:55*/;
           A_16_SS[19'h6_1ea8+7'h44] <= 16'd107;
           end 
          
      6'd55/*55:US*/:  begin 
           xpc10 <= 6'd56/*56:xpc10:56*/;
           A_16_SS[19'h6_1ea8+7'h46] <= 16'd110;
           end 
          
      6'd56/*56:US*/:  begin 
           xpc10 <= 6'd57/*57:xpc10:57*/;
           A_16_SS[19'h6_1ea8+7'h48] <= 16'd112;
           end 
          
      6'd57/*57:US*/:  begin 
           xpc10 <= 6'd58/*58:xpc10:58*/;
           A_16_SS[19'h6_1ea8+7'h4a] <= 16'd104;
           end 
          
      6'd58/*58:US*/:  begin 
           xpc10 <= 6'd59/*59:xpc10:59*/;
           A_16_SS[19'h6_1ea8+7'h4c] <= 16'd104;
           end 
          
      6'd59/*59:US*/:  begin 
           xpc10 <= 6'd60/*60:xpc10:60*/;
           A_16_SS[19'h6_1ea8+7'h4e] <= 16'd115;
           end 
          
      6'd60/*60:US*/:  begin 
           xpc10 <= 6'd61/*61:xpc10:61*/;
           A_16_SS[19'h6_1ea8+7'h50] <= 16'd113;
           end 
          
      6'd61/*61:US*/:  begin 
           xpc10 <= 6'd62/*62:xpc10:62*/;
           A_16_SS[19'h6_1ea8+7'h52] <= 16'd119;
           end 
          
      6'd62/*62:US*/:  begin 
           xpc10 <= 6'd63/*63:xpc10:63*/;
           A_16_SS[19'h6_1ea8+7'h54] <= 16'd103;
           end 
          
      6'd63/*63:US*/:  begin 
           xpc10 <= 7'd64/*64:xpc10:64*/;
           A_16_SS[19'h6_1ea8+7'h56] <= 16'd100;
           end 
          
      7'd64/*64:US*/:  begin 
           xpc10 <= 7'd65/*65:xpc10:65*/;
           A_16_SS[19'h6_1ea8+7'h58] <= 16'd109;
           end 
          
      7'd65/*65:US*/:  begin 
           xpc10 <= 7'd66/*66:xpc10:66*/;
           A_16_SS[19'h6_1ea8+7'h5a] <= 16'd107;
           end 
          
      7'd66/*66:US*/:  begin 
           xpc10 <= 7'd67/*67:xpc10:67*/;
           A_16_SS[19'h6_1ea8+7'h5c] <= 16'd108;
           end 
          
      7'd67/*67:US*/:  begin 
           xpc10 <= 7'd68/*68:xpc10:68*/;
           A_16_SS[19'h6_1ea8+7'h5e] <= 16'd121;
           end 
          
      7'd68/*68:US*/:  begin 
           xpc10 <= 7'd69/*69:xpc10:69*/;
           A_16_SS[19'h6_1ea8+7'h60] <= 16'd108;
           end 
          
      7'd69/*69:US*/:  begin 
           xpc10 <= 7'd70/*70:xpc10:70*/;
           A_16_SS[19'h6_1ea8+7'h62] <= 16'd107;
           end 
          
      7'd70/*70:US*/:  begin 
           xpc10 <= 7'd71/*71:xpc10:71*/;
           A_16_SS[19'h6_1ea8+7'h64] <= 16'd108;
           end 
          
      7'd71/*71:US*/:  begin 
           xpc10 <= 7'd72/*72:xpc10:72*/;
           A_16_SS[19'h6_1ea8+7'h66] <= 16'd113;
           end 
          
      7'd72/*72:US*/:  begin 
           xpc10 <= 7'd73/*73:xpc10:73*/;
           A_16_SS[19'h6_1ea8+7'h68] <= 16'd105;
           end 
          
      7'd73/*73:US*/:  begin 
           xpc10 <= 7'd74/*74:xpc10:74*/;
           A_16_SS[19'h6_1ea8+7'h6a] <= 16'd118;
           end 
          
      7'd74/*74:US*/:  begin 
           xpc10 <= 7'd75/*75:xpc10:75*/;
           A_16_SS[19'h6_1ea8+7'h6c] <= 16'd107;
           end 
          
      7'd75/*75:US*/:  begin 
           xpc10 <= 7'd76/*76:xpc10:76*/;
           A_16_SS[19'h6_1ea8+7'h6e] <= 16'd114;
           end 
          
      7'd76/*76:US*/:  begin 
           xpc10 <= 7'd77/*77:xpc10:77*/;
           A_16_SS[19'h6_1ea8+7'h70] <= 16'd115;
           end 
          
      7'd77/*77:US*/:  begin 
           xpc10 <= 7'd78/*78:xpc10:78*/;
           A_16_SS[19'h6_1ea8+7'h72] <= 16'd108;
           end 
          
      7'd78/*78:US*/:  begin 
           xpc10 <= 7'd79/*79:xpc10:79*/;
           A_16_SS[19'h6_1ea8+7'h74] <= 16'd101;
           end 
          
      7'd79/*79:US*/:  begin 
           xpc10 <= 7'd80/*80:xpc10:80*/;
           A_16_SS[19'h6_1ea8+7'h76] <= 16'd118;
           end 
          
      7'd80/*80:US*/:  begin 
           xpc10 <= 7'd81/*81:xpc10:81*/;
           A_16_SS[19'h6_1ea8+7'h78] <= 16'd119;
           end 
          
      7'd81/*81:US*/:  begin 
           xpc10 <= 7'd82/*82:xpc10:82*/;
           A_16_SS[19'h6_1ea8+7'h7a] <= 16'd103;
           end 
          
      7'd82/*82:US*/:  begin 
           xpc10 <= 7'd83/*83:xpc10:83*/;
           A_16_SS[19'h6_1ea8+7'h7c] <= 16'd115;
           end 
          
      7'd83/*83:US*/:  begin 
           xpc10 <= 7'd84/*84:xpc10:84*/;
           A_16_SS[19'h6_1ea8+7'h7e] <= 16'd113;
           end 
          
      7'd84/*84:US*/:  begin 
           xpc10 <= 7'd85/*85:xpc10:85*/;
           A_16_SS[19'h6_1ea8+8'h80] <= 16'd101;
           end 
          
      7'd85/*85:US*/:  begin 
           xpc10 <= 7'd86/*86:xpc10:86*/;
           A_16_SS[19'h6_1ea8+8'h82] <= 16'd97;
           end 
          
      7'd86/*86:US*/:  begin 
           xpc10 <= 7'd87/*87:xpc10:87*/;
           A_16_SS[19'h6_1ea8+8'h84] <= 16'd108;
           end 
          
      7'd87/*87:US*/:  begin 
           xpc10 <= 7'd88/*88:xpc10:88*/;
           A_16_SS[19'h6_1ea8+8'h86] <= 16'd101;
           end 
          
      7'd88/*88:US*/:  begin 
           xpc10 <= 7'd89/*89:xpc10:89*/;
           A_16_SS[19'h6_1ea8+8'h88] <= 16'd101;
           end 
          
      7'd89/*89:US*/:  begin 
           xpc10 <= 7'd90/*90:xpc10:90*/;
           A_16_SS[19'h6_1ea8+8'h8a] <= 16'd97;
           end 
          
      7'd90/*90:US*/:  begin 
           xpc10 <= 7'd91/*91:xpc10:91*/;
           A_16_SS[19'h6_1ea8+8'h8c] <= 16'd107;
           end 
          
      7'd91/*91:US*/:  begin 
           xpc10 <= 7'd92/*92:xpc10:92*/;
           A_16_SS[19'h6_1ea8+8'h8e] <= 16'd101;
           end 
          
      7'd92/*92:US*/:  begin 
           xpc10 <= 7'd93/*93:xpc10:93*/;
           A_16_SS[19'h6_1ea8+8'h90] <= 16'd118;
           end 
          
      7'd93/*93:US*/:  begin 
           xpc10 <= 7'd94/*94:xpc10:94*/;
           A_16_SS[19'h6_1ea8+8'h92] <= 16'd114;
           end 
          
      7'd94/*94:US*/:  begin 
           xpc10 <= 7'd95/*95:xpc10:95*/;
           A_16_SS[19'h6_1ea8+8'h94] <= 16'd113;
           end 
          
      7'd95/*95:US*/:  begin 
           xpc10 <= 7'd96/*96:xpc10:96*/;
           A_16_SS[19'h6_1ea8+8'h96] <= 16'd101;
           end 
          
      7'd96/*96:US*/:  begin 
           xpc10 <= 7'd97/*97:xpc10:97*/;
           A_16_SS[19'h6_1ea8+8'h98] <= 16'd110;
           end 
          
      7'd97/*97:US*/:  begin 
           xpc10 <= 7'd98/*98:xpc10:98*/;
           A_16_SS[19'h6_1f42+0] <= 16'd112;
           end 
          
      7'd98/*98:US*/:  begin 
           xpc10 <= 7'd99/*99:xpc10:99*/;
           A_16_SS[19'h6_1f42+2'h2] <= 16'd112;
           end 
          
      7'd99/*99:US*/:  begin 
           xpc10 <= 7'd100/*100:xpc10:100*/;
           A_16_SS[19'h6_1f42+3'h4] <= 16'd101;
           end 
          
      7'd100/*100:US*/:  begin 
           xpc10 <= 7'd101/*101:xpc10:101*/;
           A_16_SS[19'h6_1f42+3'h6] <= 16'd97;
           end 
          
      7'd101/*101:US*/:  begin 
           xpc10 <= 7'd102/*102:xpc10:102*/;
           A_16_SS[19'h6_1f42+4'h8] <= 16'd105;
           end 
          
      7'd102/*102:US*/:  begin 
           xpc10 <= 7'd103/*103:xpc10:103*/;
           A_16_SS[19'h6_1f42+4'ha] <= 16'd112;
           end 
          
      7'd103/*103:US*/:  begin 
           xpc10 <= 7'd104/*104:xpc10:104*/;
           A_16_SS[19'h6_1f42+4'hc] <= 16'd102;
           end 
          
      7'd104/*104:US*/:  begin 
           xpc10 <= 7'd105/*105:xpc10:105*/;
           A_16_SS[19'h6_1f42+4'he] <= 16'd114;
           end 
          
      7'd105/*105:US*/:  begin 
           xpc10 <= 7'd106/*106:xpc10:106*/;
           A_16_SS[19'h6_1f42+5'h10] <= 16'd112;
           end 
          
      7'd106/*106:US*/:  begin 
           xpc10 <= 7'd107/*107:xpc10:107*/;
           A_16_SS[19'h6_1f42+5'h12] <= 16'd101;
           end 
          
      7'd107/*107:US*/:  begin 
           xpc10 <= 7'd108/*108:xpc10:108*/;
           A_16_SS[19'h6_1f42+5'h14] <= 16'd121;
           end 
          
      7'd108/*108:US*/:  begin 
           xpc10 <= 7'd109/*109:xpc10:109*/;
           A_16_SS[19'h6_1f42+5'h16] <= 16'd97;
           end 
          
      7'd109/*109:US*/:  begin 
           xpc10 <= 7'd110/*110:xpc10:110*/;
           A_16_SS[19'h6_1f42+5'h18] <= 16'd110;
           end 
          
      7'd110/*110:US*/:  begin 
           xpc10 <= 7'd111/*111:xpc10:111*/;
           A_16_SS[19'h6_1f42+5'h1a] <= 16'd114;
           end 
          
      7'd111/*111:US*/:  begin 
           xpc10 <= 7'd112/*112:xpc10:112*/;
           A_16_SS[19'h6_1f42+5'h1c] <= 16'd108;
           end 
          
      7'd112/*112:US*/:  begin 
           xpc10 <= 7'd113/*113:xpc10:113*/;
           A_16_SS[19'h6_1f42+5'h1e] <= 16'd108;
           end 
          
      7'd113/*113:US*/:  begin 
           xpc10 <= 7'd114/*114:xpc10:114*/;
           A_16_SS[19'h6_1f42+6'h20] <= 16'd103;
           end 
          
      7'd114/*114:US*/:  begin 
           xpc10 <= 7'd115/*115:xpc10:115*/;
           A_16_SS[19'h6_1f42+6'h22] <= 16'd116;
           end 
          
      7'd115/*115:US*/:  begin 
           xpc10 <= 7'd116/*116:xpc10:116*/;
           A_16_SS[19'h6_1f42+6'h24] <= 16'd115;
           end 
          
      7'd116/*116:US*/:  begin 
           xpc10 <= 7'd117/*117:xpc10:117*/;
           A_16_SS[19'h6_1f42+6'h26] <= 16'd121;
           end 
          
      7'd117/*117:US*/:  begin 
           xpc10 <= 7'd118/*118:xpc10:118*/;
           A_16_SS[19'h6_1f42+6'h28] <= 16'd112;
           end 
          
      7'd118/*118:US*/:  begin 
           xpc10 <= 7'd119/*119:xpc10:119*/;
           A_16_SS[19'h6_1f42+6'h2a] <= 16'd101;
           end 
          
      7'd119/*119:US*/:  begin 
           xpc10 <= 7'd120/*120:xpc10:120*/;
           A_16_SS[19'h6_1f42+6'h2c] <= 16'd97;
           end 
          
      7'd120/*120:US*/:  begin 
           xpc10 <= 7'd121/*121:xpc10:121*/;
           A_16_SS[19'h6_1f42+6'h2e] <= 16'd101;
           end 
          
      7'd121/*121:US*/:  begin 
           xpc10 <= 7'd122/*122:xpc10:122*/;
           A_16_SS[19'h6_1f42+6'h30] <= 16'd113;
           end 
          
      7'd122/*122:US*/:  begin 
           xpc10 <= 7'd123/*123:xpc10:123*/;
           A_16_SS[19'h6_1f42+6'h32] <= 16'd105;
           end 
          
      7'd123/*123:US*/:  begin 
           xpc10 <= 7'd124/*124:xpc10:124*/;
           A_16_SS[19'h6_1f42+6'h34] <= 16'd97;
           end 
          
      7'd124/*124:US*/:  begin 
           xpc10 <= 7'd125/*125:xpc10:125*/;
           A_16_SS[19'h6_1f42+6'h36] <= 16'd105;
           end 
          
      7'd125/*125:US*/:  begin 
           xpc10 <= 7'd126/*126:xpc10:126*/;
           A_16_SS[19'h6_1f42+6'h38] <= 16'd108;
           end 
          
      7'd126/*126:US*/:  begin 
           xpc10 <= 7'd127/*127:xpc10:127*/;
           A_16_SS[19'h6_1f42+6'h3a] <= 16'd107;
           end 
          
      7'd127/*127:US*/:  begin 
           xpc10 <= 8'd128/*128:xpc10:128*/;
           A_16_SS[19'h6_1f42+6'h3c] <= 16'd114;
           end 
          
      8'd128/*128:US*/:  begin 
           xpc10 <= 8'd129/*129:xpc10:129*/;
           A_16_SS[19'h6_1f42+6'h3e] <= 16'd108;
           end 
          
      8'd129/*129:US*/:  begin 
           xpc10 <= 8'd130/*130:xpc10:130*/;
           A_16_SS[19'h6_1f42+7'h40] <= 16'd103;
           end 
          
      8'd130/*130:US*/:  begin 
           xpc10 <= 8'd131/*131:xpc10:131*/;
           A_16_SS[19'h6_1f42+7'h42] <= 16'd99;
           end 
          
      8'd131/*131:US*/:  begin 
           xpc10 <= 8'd132/*132:xpc10:132*/;
           A_16_SS[19'h6_1f42+7'h44] <= 16'd114;
           end 
          
      8'd132/*132:US*/:  begin 
           xpc10 <= 8'd133/*133:xpc10:133*/;
           A_16_SS[19'h6_1f42+7'h46] <= 16'd118;
           end 
          
      8'd133/*133:US*/:  begin 
           xpc10 <= 8'd134/*134:xpc10:134*/;
           A_16_SS[19'h6_1f42+7'h48] <= 16'd101;
           end 
          
      8'd134/*134:US*/:  begin 
           xpc10 <= 8'd135/*135:xpc10:135*/;
           A_16_SS[19'h6_1f42+7'h4a] <= 16'd103;
           end 
          
      8'd135/*135:US*/:  begin 
           xpc10 <= 8'd136/*136:xpc10:136*/;
           A_16_SS[19'h6_1f42+7'h4c] <= 16'd101;
           end 
          
      8'd136/*136:US*/:  begin 
           xpc10 <= 8'd137/*137:xpc10:137*/;
           A_16_SS[19'h6_1f42+7'h4e] <= 16'd103;
           end 
          
      8'd137/*137:US*/:  begin 
           xpc10 <= 8'd138/*138:xpc10:138*/;
           A_16_SS[19'h6_1f42+7'h50] <= 16'd112;
           end 
          
      8'd138/*138:US*/:  begin 
           xpc10 <= 8'd139/*139:xpc10:139*/;
           A_16_SS[19'h6_1f42+7'h52] <= 16'd116;
           end 
          
      8'd139/*139:US*/:  begin 
           xpc10 <= 8'd140/*140:xpc10:140*/;
           A_16_SS[19'h6_1f42+7'h54] <= 16'd121;
           end 
          
      8'd140/*140:US*/:  begin 
           xpc10 <= 8'd141/*141:xpc10:141*/;
           A_16_SS[19'h6_1f42+7'h56] <= 16'd114;
           end 
          
      8'd141/*141:US*/:  begin 
           xpc10 <= 8'd142/*142:xpc10:142*/;
           A_16_SS[19'h6_1f42+7'h58] <= 16'd118;
           end 
          
      8'd142/*142:US*/:  begin 
           xpc10 <= 8'd143/*143:xpc10:143*/;
           A_16_SS[19'h6_1f42+7'h5a] <= 16'd116;
           end 
          
      8'd143/*143:US*/:  begin 
           xpc10 <= 8'd144/*144:xpc10:144*/;
           A_16_SS[19'h6_1f42+7'h5c] <= 16'd112;
           end 
          
      8'd144/*144:US*/:  begin 
           xpc10 <= 8'd145/*145:xpc10:145*/;
           A_16_SS[19'h6_1f42+7'h5e] <= 16'd112;
           end 
          
      8'd145/*145:US*/:  begin 
           xpc10 <= 8'd146/*146:xpc10:146*/;
           A_16_SS[19'h6_1f42+7'h60] <= 16'd115;
           end 
          
      8'd146/*146:US*/:  begin 
           xpc10 <= 8'd147/*147:xpc10:147*/;
           A_16_SS[19'h6_1f42+7'h62] <= 16'd104;
           end 
          
      8'd147/*147:US*/:  begin 
           xpc10 <= 8'd148/*148:xpc10:148*/;
           A_16_SS[19'h6_1f42+7'h64] <= 16'd114;
           end 
          
      8'd148/*148:US*/:  begin 
           xpc10 <= 8'd149/*149:xpc10:149*/;
           A_16_SS[19'h6_1f42+7'h66] <= 16'd108;
           end 
          
      8'd149/*149:US*/:  begin 
           xpc10 <= 8'd150/*150:xpc10:150*/;
           A_16_SS[19'h6_1f42+7'h68] <= 16'd100;
           end 
          
      8'd150/*150:US*/:  begin 
           xpc10 <= 8'd151/*151:xpc10:151*/;
           A_16_SS[19'h6_1f42+7'h6a] <= 16'd108;
           end 
          
      8'd151/*151:US*/:  begin 
           xpc10 <= 8'd152/*152:xpc10:152*/;
           A_16_SS[19'h6_1f42+7'h6c] <= 16'd114;
           end 
          
      8'd152/*152:US*/:  begin 
           xpc10 <= 8'd153/*153:xpc10:153*/;
           A_16_SS[19'h6_1f42+7'h6e] <= 16'd108;
           end 
          
      8'd153/*153:US*/:  begin 
           xpc10 <= 8'd154/*154:xpc10:154*/;
           A_16_SS[19'h6_1f42+7'h70] <= 16'd101;
           end 
          
      8'd154/*154:US*/:  begin 
           xpc10 <= 8'd155/*155:xpc10:155*/;
           A_16_SS[19'h6_1f42+7'h72] <= 16'd101;
           end 
          
      8'd155/*155:US*/:  begin 
           xpc10 <= 8'd156/*156:xpc10:156*/;
           A_16_SS[19'h6_1f42+7'h74] <= 16'd100;
           end 
          
      8'd156/*156:US*/:  begin 
           xpc10 <= 8'd157/*157:xpc10:157*/;
           A_16_SS[19'h6_1f42+7'h76] <= 16'd108;
           end 
          
      8'd157/*157:US*/:  begin 
           xpc10 <= 8'd158/*158:xpc10:158*/;
           A_16_SS[19'h6_1f42+7'h78] <= 16'd118;
           end 
          
      8'd158/*158:US*/:  begin 
           xpc10 <= 8'd159/*159:xpc10:159*/;
           A_16_SS[19'h6_1f42+7'h7a] <= 16'd101;
           end 
          
      8'd159/*159:US*/:  begin 
           xpc10 <= 8'd160/*160:xpc10:160*/;
           A_16_SS[19'h6_1f42+7'h7c] <= 16'd101;
           end 
          
      8'd160/*160:US*/:  begin 
           xpc10 <= 8'd161/*161:xpc10:161*/;
           A_16_SS[19'h6_1f42+7'h7e] <= 16'd118;
           end 
          
      8'd161/*161:US*/:  begin 
           xpc10 <= 8'd162/*162:xpc10:162*/;
           A_16_SS[19'h6_1f42+8'h80] <= 16'd97;
           end 
          
      8'd162/*162:US*/:  begin 
           xpc10 <= 8'd163/*163:xpc10:163*/;
           A_16_SS[19'h6_1f42+8'h82] <= 16'd114;
           end 
          
      8'd163/*163:US*/:  begin 
           xpc10 <= 8'd164/*164:xpc10:164*/;
           A_16_SS[19'h6_1f42+8'h84] <= 16'd105;
           end 
          
      8'd164/*164:US*/:  begin 
           xpc10 <= 8'd165/*165:xpc10:165*/;
           A_16_SS[19'h6_1f42+8'h86] <= 16'd113;
           end 
          
      8'd165/*165:US*/:  begin 
           xpc10 <= 8'd166/*166:xpc10:166*/;
           A_16_SS[19'h6_1f42+8'h88] <= 16'd103;
           end 
          
      8'd166/*166:US*/:  begin 
           xpc10 <= 8'd167/*167:xpc10:167*/;
           A_16_SS[19'h6_1f42+8'h8a] <= 16'd121;
           end 
          
      8'd167/*167:US*/:  begin 
           xpc10 <= 8'd168/*168:xpc10:168*/;
           A_16_SS[19'h6_1f42+8'h8c] <= 16'd101;
           end 
          
      8'd168/*168:US*/:  begin 
           xpc10 <= 8'd169/*169:xpc10:169*/;
           A_16_SS[19'h6_1f42+8'h8e] <= 16'd116;
           end 
          
      8'd169/*169:US*/:  begin 
           xpc10 <= 8'd170/*170:xpc10:170*/;
           A_16_SS[19'h6_1f42+8'h90] <= 16'd105;
           end 
          
      8'd170/*170:US*/:  begin 
           xpc10 <= 8'd171/*171:xpc10:171*/;
           A_16_SS[19'h6_1f42+8'h92] <= 16'd112;
           end 
          
      8'd171/*171:US*/:  begin 
           xpc10 <= 8'd172/*172:xpc10:172*/;
           A_SINT[64'h6_1fd8+64'd4] <= 32'd20;
           A_16_SS[19'h6_1f42+8'h94] <= 16'd108;
           end 
          
      8'd172/*172:US*/:  begin 
           xpc10 <= 8'd173/*173:xpc10:173*/;
           A_SINT[19'h6_1fd8+4'd8] <= 32'd20;
           end 
          
      8'd173/*173:US*/:  begin 
           xpc10 <= 8'd174/*174:xpc10:174*/;
           A_SINT[19'h6_1fe8+0] <= 32'd2;
           end 
          
      8'd174/*174:US*/:  begin 
           xpc10 <= 8'd175/*175:xpc10:175*/;
           A_SINT[19'h6_1fe8+3'h4] <= -32'd2;
           end 
          
      8'd175/*175:US*/:  begin 
           xpc10 <= 8'd176/*176:xpc10:176*/;
           A_SINT[19'h6_1fe8+4'h8] <= 32'd0;
           end 
          
      8'd176/*176:US*/:  begin 
           xpc10 <= 8'd177/*177:xpc10:177*/;
           A_SINT[19'h6_1fe8+4'hc] <= 32'd0;
           end 
          
      8'd177/*177:US*/:  begin 
           xpc10 <= 8'd178/*178:xpc10:178*/;
           A_SINT[19'h6_1fe8+5'h10] <= -32'd4;
           end 
          
      8'd178/*178:US*/:  begin 
           xpc10 <= 8'd179/*179:xpc10:179*/;
           A_SINT[19'h6_1fe8+5'h14] <= 32'd1;
           end 
          
      8'd179/*179:US*/:  begin 
           xpc10 <= 8'd180/*180:xpc10:180*/;
           A_SINT[19'h6_1fe8+5'h18] <= -32'd1;
           end 
          
      8'd180/*180:US*/:  begin 
           xpc10 <= 8'd181/*181:xpc10:181*/;
           A_SINT[19'h6_1fe8+5'h1c] <= -32'd1;
           end 
          
      8'd181/*181:US*/:  begin 
           xpc10 <= 8'd182/*182:xpc10:182*/;
           A_SINT[19'h6_1fe8+6'h20] <= -32'd1;
           end 
          
      8'd182/*182:US*/:  begin 
           xpc10 <= 8'd183/*183:xpc10:183*/;
           A_SINT[19'h6_1fe8+6'h24] <= -32'd2;
           end 
          
      8'd183/*183:US*/:  begin 
           xpc10 <= 8'd184/*184:xpc10:184*/;
           A_SINT[19'h6_1fe8+6'h28] <= -32'd1;
           end 
          
      8'd184/*184:US*/:  begin 
           xpc10 <= 8'd185/*185:xpc10:185*/;
           A_SINT[19'h6_1fe8+6'h2c] <= 32'd0;
           end 
          
      8'd185/*185:US*/:  begin 
           xpc10 <= 8'd186/*186:xpc10:186*/;
           A_SINT[19'h6_1fe8+6'h30] <= 32'd1;
           end 
          
      8'd186/*186:US*/:  begin 
           xpc10 <= 8'd187/*187:xpc10:187*/;
           A_SINT[19'h6_1fe8+6'h34] <= 32'd0;
           end 
          
      8'd187/*187:US*/:  begin 
           xpc10 <= 8'd188/*188:xpc10:188*/;
           A_SINT[19'h6_1fe8+6'h38] <= -32'd2;
           end 
          
      8'd188/*188:US*/:  begin 
           xpc10 <= 8'd189/*189:xpc10:189*/;
           A_SINT[19'h6_1fe8+6'h3c] <= 32'd1;
           end 
          
      8'd189/*189:US*/:  begin 
           xpc10 <= 8'd190/*190:xpc10:190*/;
           A_SINT[19'h6_1fe8+7'h40] <= 32'd1;
           end 
          
      8'd190/*190:US*/:  begin 
           xpc10 <= 8'd191/*191:xpc10:191*/;
           A_SINT[19'h6_1fe8+7'h44] <= 32'd0;
           end 
          
      8'd191/*191:US*/:  begin 
           xpc10 <= 8'd192/*192:xpc10:192*/;
           A_SINT[19'h6_1fe8+7'h48] <= -32'd1;
           end 
          
      8'd192/*192:US*/:  begin 
           xpc10 <= 8'd193/*193:xpc10:193*/;
           A_SINT[19'h6_1fe8+7'h4c] <= -32'd3;
           end 
          
      8'd193/*193:US*/:  begin 
           xpc10 <= 8'd194/*194:xpc10:194*/;
           A_SINT[19'h6_1fe8+7'h50] <= -32'd2;
           end 
          
      8'd194/*194:US*/:  begin 
           xpc10 <= 8'd195/*195:xpc10:195*/;
           A_SINT[19'h6_1fe8+7'h54] <= 32'd12;
           end 
          
      8'd195/*195:US*/:  begin 
           xpc10 <= 8'd196/*196:xpc10:196*/;
           A_SINT[19'h6_1fe8+7'h58] <= -32'd5;
           end 
          
      8'd196/*196:US*/:  begin 
           xpc10 <= 8'd197/*197:xpc10:197*/;
           A_SINT[19'h6_1fe8+7'h5c] <= -32'd5;
           end 
          
      8'd197/*197:US*/:  begin 
           xpc10 <= 8'd198/*198:xpc10:198*/;
           A_SINT[19'h6_1fe8+7'h60] <= -32'd4;
           end 
          
      8'd198/*198:US*/:  begin 
           xpc10 <= 8'd199/*199:xpc10:199*/;
           A_SINT[19'h6_1fe8+7'h64] <= -32'd3;
           end 
          
      8'd199/*199:US*/:  begin 
           xpc10 <= 8'd200/*200:xpc10:200*/;
           A_SINT[19'h6_1fe8+7'h68] <= -32'd3;
           end 
          
      8'd200/*200:US*/:  begin 
           xpc10 <= 8'd201/*201:xpc10:201*/;
           A_SINT[19'h6_1fe8+7'h6c] <= -32'd2;
           end 
          
      8'd201/*201:US*/:  begin 
           xpc10 <= 8'd202/*202:xpc10:202*/;
           A_SINT[19'h6_1fe8+7'h70] <= -32'd5;
           end 
          
      8'd202/*202:US*/:  begin 
           xpc10 <= 8'd203/*203:xpc10:203*/;
           A_SINT[19'h6_1fe8+7'h74] <= -32'd6;
           end 
          
      8'd203/*203:US*/:  begin 
           xpc10 <= 8'd204/*204:xpc10:204*/;
           A_SINT[19'h6_1fe8+7'h78] <= -32'd5;
           end 
          
      8'd204/*204:US*/:  begin 
           xpc10 <= 8'd205/*205:xpc10:205*/;
           A_SINT[19'h6_1fe8+7'h7c] <= -32'd4;
           end 
          
      8'd205/*205:US*/:  begin 
           xpc10 <= 8'd206/*206:xpc10:206*/;
           A_SINT[19'h6_1fe8+8'h80] <= -32'd3;
           end 
          
      8'd206/*206:US*/:  begin 
           xpc10 <= 8'd207/*207:xpc10:207*/;
           A_SINT[19'h6_1fe8+8'h84] <= -32'd5;
           end 
          
      8'd207/*207:US*/:  begin 
           xpc10 <= 8'd208/*208:xpc10:208*/;
           A_SINT[19'h6_1fe8+8'h88] <= -32'd4;
           end 
          
      8'd208/*208:US*/:  begin 
           xpc10 <= 8'd209/*209:xpc10:209*/;
           A_SINT[19'h6_1fe8+8'h8c] <= 32'd0;
           end 
          
      8'd209/*209:US*/:  begin 
           xpc10 <= 8'd210/*210:xpc10:210*/;
           A_SINT[19'h6_1fe8+8'h90] <= -32'd2;
           end 
          
      8'd210/*210:US*/:  begin 
           xpc10 <= 8'd211/*211:xpc10:211*/;
           A_SINT[19'h6_1fe8+8'h94] <= -32'd2;
           end 
          
      8'd211/*211:US*/:  begin 
           xpc10 <= 8'd212/*212:xpc10:212*/;
           A_SINT[19'h6_1fe8+8'h98] <= -32'd8;
           end 
          
      8'd212/*212:US*/:  begin 
           xpc10 <= 8'd213/*213:xpc10:213*/;
           A_SINT[19'h6_1fe8+8'h9c] <= 32'd0;
           end 
          
      8'd213/*213:US*/:  begin 
           xpc10 <= 8'd214/*214:xpc10:214*/;
           A_SINT[19'h6_1fe8+8'ha0] <= 32'd0;
           end 
          
      8'd214/*214:US*/:  begin 
           xpc10 <= 8'd215/*215:xpc10:215*/;
           A_SINT[19'h6_1fe8+8'ha4] <= -32'd5;
           end 
          
      8'd215/*215:US*/:  begin 
           xpc10 <= 8'd216/*216:xpc10:216*/;
           A_SINT[19'h6_1fe8+8'ha8] <= 32'd4;
           end 
          
      8'd216/*216:US*/:  begin 
           xpc10 <= 8'd217/*217:xpc10:217*/;
           A_SINT[19'h6_1fe8+8'hac] <= 32'd3;
           end 
          
      8'd217/*217:US*/:  begin 
           xpc10 <= 8'd218/*218:xpc10:218*/;
           A_SINT[19'h6_1fe8+8'hb0] <= -32'd6;
           end 
          
      8'd218/*218:US*/:  begin 
           xpc10 <= 8'd219/*219:xpc10:219*/;
           A_SINT[19'h6_1fe8+8'hb4] <= 32'd1;
           end 
          
      8'd219/*219:US*/:  begin 
           xpc10 <= 8'd220/*220:xpc10:220*/;
           A_SINT[19'h6_1fe8+8'hb8] <= 32'd1;
           end 
          
      8'd220/*220:US*/:  begin 
           xpc10 <= 8'd221/*221:xpc10:221*/;
           A_SINT[19'h6_1fe8+8'hbc] <= -32'd2;
           end 
          
      8'd221/*221:US*/:  begin 
           xpc10 <= 8'd222/*222:xpc10:222*/;
           A_SINT[19'h6_1fe8+8'hc0] <= 32'd0;
           end 
          
      8'd222/*222:US*/:  begin 
           xpc10 <= 8'd223/*223:xpc10:223*/;
           A_SINT[19'h6_1fe8+8'hc4] <= -32'd4;
           end 
          
      8'd223/*223:US*/:  begin 
           xpc10 <= 8'd224/*224:xpc10:224*/;
           A_SINT[19'h6_1fe8+8'hc8] <= -32'd3;
           end 
          
      8'd224/*224:US*/:  begin 
           xpc10 <= 8'd225/*225:xpc10:225*/;
           A_SINT[19'h6_1fe8+8'hcc] <= 32'd2;
           end 
          
      8'd225/*225:US*/:  begin 
           xpc10 <= 8'd226/*226:xpc10:226*/;
           A_SINT[19'h6_1fe8+8'hd0] <= -32'd1;
           end 
          
      8'd226/*226:US*/:  begin 
           xpc10 <= 8'd227/*227:xpc10:227*/;
           A_SINT[19'h6_1fe8+8'hd4] <= 32'd2;
           end 
          
      8'd227/*227:US*/:  begin 
           xpc10 <= 8'd228/*228:xpc10:228*/;
           A_SINT[19'h6_1fe8+8'hd8] <= -32'd1;
           end 
          
      8'd228/*228:US*/:  begin 
           xpc10 <= 8'd229/*229:xpc10:229*/;
           A_SINT[19'h6_1fe8+8'hdc] <= 32'd0;
           end 
          
      8'd229/*229:US*/:  begin 
           xpc10 <= 8'd230/*230:xpc10:230*/;
           A_SINT[19'h6_1fe8+8'he0] <= 32'd0;
           end 
          
      8'd230/*230:US*/:  begin 
           xpc10 <= 8'd231/*231:xpc10:231*/;
           A_SINT[19'h6_1fe8+8'he4] <= -32'd2;
           end 
          
      8'd231/*231:US*/:  begin 
           xpc10 <= 8'd232/*232:xpc10:232*/;
           A_SINT[19'h6_1fe8+8'he8] <= -32'd7;
           end 
          
      8'd232/*232:US*/:  begin 
           xpc10 <= 8'd233/*233:xpc10:233*/;
           A_SINT[19'h6_1fe8+8'hec] <= -32'd4;
           end 
          
      8'd233/*233:US*/:  begin 
           xpc10 <= 8'd234/*234:xpc10:234*/;
           A_SINT[19'h6_1fe8+8'hf0] <= 32'd0;
           end 
          
      8'd234/*234:US*/:  begin 
           xpc10 <= 8'd235/*235:xpc10:235*/;
           A_SINT[19'h6_1fe8+8'hf4] <= -32'd5;
           end 
          
      8'd235/*235:US*/:  begin 
           xpc10 <= 8'd236/*236:xpc10:236*/;
           A_SINT[19'h6_1fe8+8'hf8] <= 32'd3;
           end 
          
      8'd236/*236:US*/:  begin 
           xpc10 <= 8'd237/*237:xpc10:237*/;
           A_SINT[19'h6_1fe8+8'hfc] <= 32'd4;
           end 
          
      8'd237/*237:US*/:  begin 
           xpc10 <= 8'd238/*238:xpc10:238*/;
           A_SINT[19'h6_1fe8+9'h100] <= -32'd5;
           end 
          
      8'd238/*238:US*/:  begin 
           xpc10 <= 8'd239/*239:xpc10:239*/;
           A_SINT[19'h6_1fe8+9'h104] <= 32'd0;
           end 
          
      8'd239/*239:US*/:  begin 
           xpc10 <= 8'd240/*240:xpc10:240*/;
           A_SINT[19'h6_1fe8+9'h108] <= 32'd1;
           end 
          
      8'd240/*240:US*/:  begin 
           xpc10 <= 8'd241/*241:xpc10:241*/;
           A_SINT[19'h6_1fe8+9'h10c] <= -32'd2;
           end 
          
      8'd241/*241:US*/:  begin 
           xpc10 <= 8'd242/*242:xpc10:242*/;
           A_SINT[19'h6_1fe8+9'h110] <= 32'd0;
           end 
          
      8'd242/*242:US*/:  begin 
           xpc10 <= 8'd243/*243:xpc10:243*/;
           A_SINT[19'h6_1fe8+9'h114] <= -32'd3;
           end 
          
      8'd243/*243:US*/:  begin 
           xpc10 <= 8'd244/*244:xpc10:244*/;
           A_SINT[19'h6_1fe8+9'h118] <= -32'd2;
           end 
          
      8'd244/*244:US*/:  begin 
           xpc10 <= 8'd245/*245:xpc10:245*/;
           A_SINT[19'h6_1fe8+9'h11c] <= 32'd1;
           end 
          
      8'd245/*245:US*/:  begin 
           xpc10 <= 8'd246/*246:xpc10:246*/;
           A_SINT[19'h6_1fe8+9'h120] <= -32'd1;
           end 
          
      8'd246/*246:US*/:  begin 
           xpc10 <= 8'd247/*247:xpc10:247*/;
           A_SINT[19'h6_1fe8+9'h124] <= 32'd2;
           end 
          
      8'd247/*247:US*/:  begin 
           xpc10 <= 8'd248/*248:xpc10:248*/;
           A_SINT[19'h6_1fe8+9'h128] <= -32'd1;
           end 
          
      8'd248/*248:US*/:  begin 
           xpc10 <= 8'd249/*249:xpc10:249*/;
           A_SINT[19'h6_1fe8+9'h12c] <= 32'd0;
           end 
          
      8'd249/*249:US*/:  begin 
           xpc10 <= 8'd250/*250:xpc10:250*/;
           A_SINT[19'h6_1fe8+9'h130] <= 32'd0;
           end 
          
      8'd250/*250:US*/:  begin 
           xpc10 <= 8'd251/*251:xpc10:251*/;
           A_SINT[19'h6_1fe8+9'h134] <= -32'd2;
           end 
          
      8'd251/*251:US*/:  begin 
           xpc10 <= 8'd252/*252:xpc10:252*/;
           A_SINT[19'h6_1fe8+9'h138] <= -32'd7;
           end 
          
      8'd252/*252:US*/:  begin 
           xpc10 <= 8'd253/*253:xpc10:253*/;
           A_SINT[19'h6_1fe8+9'h13c] <= -32'd4;
           end 
          
      8'd253/*253:US*/:  begin 
           xpc10 <= 8'd254/*254:xpc10:254*/;
           A_SINT[19'h6_1fe8+9'h140] <= -32'd4;
           end 
          
      8'd254/*254:US*/:  begin 
           xpc10 <= 8'd255/*255:xpc10:255*/;
           A_SINT[19'h6_1fe8+9'h144] <= -32'd4;
           end 
          
      8'd255/*255:US*/:  begin 
           xpc10 <= 9'd256/*256:xpc10:256*/;
           A_SINT[19'h6_1fe8+9'h148] <= -32'd6;
           end 
          
      9'd256/*256:US*/:  begin 
           xpc10 <= 9'd257/*257:xpc10:257*/;
           A_SINT[19'h6_1fe8+9'h14c] <= -32'd5;
           end 
          
      9'd257/*257:US*/:  begin 
           xpc10 <= 9'd258/*258:xpc10:258*/;
           A_SINT[19'h6_1fe8+9'h150] <= 32'd9;
           end 
          
      9'd258/*258:US*/:  begin 
           xpc10 <= 9'd259/*259:xpc10:259*/;
           A_SINT[19'h6_1fe8+9'h154] <= -32'd5;
           end 
          
      9'd259/*259:US*/:  begin 
           xpc10 <= 9'd260/*260:xpc10:260*/;
           A_SINT[19'h6_1fe8+9'h158] <= -32'd2;
           end 
          
      9'd260/*260:US*/:  begin 
           xpc10 <= 9'd261/*261:xpc10:261*/;
           A_SINT[19'h6_1fe8+9'h15c] <= 32'd1;
           end 
          
      9'd261/*261:US*/:  begin 
           xpc10 <= 9'd262/*262:xpc10:262*/;
           A_SINT[19'h6_1fe8+9'h160] <= -32'd5;
           end 
          
      9'd262/*262:US*/:  begin 
           xpc10 <= 9'd263/*263:xpc10:263*/;
           A_SINT[19'h6_1fe8+9'h164] <= 32'd2;
           end 
          
      9'd263/*263:US*/:  begin 
           xpc10 <= 9'd264/*264:xpc10:264*/;
           A_SINT[19'h6_1fe8+9'h168] <= 32'd0;
           end 
          
      9'd264/*264:US*/:  begin 
           xpc10 <= 9'd265/*265:xpc10:265*/;
           A_SINT[19'h6_1fe8+9'h16c] <= -32'd4;
           end 
          
      9'd265/*265:US*/:  begin 
           xpc10 <= 9'd266/*266:xpc10:266*/;
           A_SINT[19'h6_1fe8+9'h170] <= -32'd5;
           end 
          
      9'd266/*266:US*/:  begin 
           xpc10 <= 9'd267/*267:xpc10:267*/;
           A_SINT[19'h6_1fe8+9'h174] <= -32'd5;
           end 
          
      9'd267/*267:US*/:  begin 
           xpc10 <= 9'd268/*268:xpc10:268*/;
           A_SINT[19'h6_1fe8+9'h178] <= -32'd4;
           end 
          
      9'd268/*268:US*/:  begin 
           xpc10 <= 9'd269/*269:xpc10:269*/;
           A_SINT[19'h6_1fe8+9'h17c] <= -32'd3;
           end 
          
      9'd269/*269:US*/:  begin 
           xpc10 <= 9'd270/*270:xpc10:270*/;
           A_SINT[19'h6_1fe8+9'h180] <= -32'd3;
           end 
          
      9'd270/*270:US*/:  begin 
           xpc10 <= 9'd271/*271:xpc10:271*/;
           A_SINT[19'h6_1fe8+9'h184] <= -32'd1;
           end 
          
      9'd271/*271:US*/:  begin 
           xpc10 <= 9'd272/*272:xpc10:272*/;
           A_SINT[19'h6_1fe8+9'h188] <= 32'd0;
           end 
          
      9'd272/*272:US*/:  begin 
           xpc10 <= 9'd273/*273:xpc10:273*/;
           A_SINT[19'h6_1fe8+9'h18c] <= 32'd7;
           end 
          
      9'd273/*273:US*/:  begin 
           xpc10 <= 9'd274/*274:xpc10:274*/;
           A_SINT[19'h6_1fe8+9'h190] <= 32'd1;
           end 
          
      9'd274/*274:US*/:  begin 
           xpc10 <= 9'd275/*275:xpc10:275*/;
           A_SINT[19'h6_1fe8+9'h194] <= -32'd3;
           end 
          
      9'd275/*275:US*/:  begin 
           xpc10 <= 9'd276/*276:xpc10:276*/;
           A_SINT[19'h6_1fe8+9'h198] <= 32'd1;
           end 
          
      9'd276/*276:US*/:  begin 
           xpc10 <= 9'd277/*277:xpc10:277*/;
           A_SINT[19'h6_1fe8+9'h19c] <= 32'd0;
           end 
          
      9'd277/*277:US*/:  begin 
           xpc10 <= 9'd278/*278:xpc10:278*/;
           A_SINT[19'h6_1fe8+9'h1a0] <= -32'd5;
           end 
          
      9'd278/*278:US*/:  begin 
           xpc10 <= 9'd279/*279:xpc10:279*/;
           A_SINT[19'h6_1fe8+9'h1a4] <= 32'd5;
           end 
          
      9'd279/*279:US*/:  begin 
           xpc10 <= 9'd280/*280:xpc10:280*/;
           A_SINT[19'h6_1fe8+9'h1a8] <= -32'd2;
           end 
          
      9'd280/*280:US*/:  begin 
           xpc10 <= 9'd281/*281:xpc10:281*/;
           A_SINT[19'h6_1fe8+9'h1ac] <= -32'd3;
           end 
          
      9'd281/*281:US*/:  begin 
           xpc10 <= 9'd282/*282:xpc10:282*/;
           A_SINT[19'h6_1fe8+9'h1b0] <= -32'd2;
           end 
          
      9'd282/*282:US*/:  begin 
           xpc10 <= 9'd283/*283:xpc10:283*/;
           A_SINT[19'h6_1fe8+9'h1b4] <= -32'd4;
           end 
          
      9'd283/*283:US*/:  begin 
           xpc10 <= 9'd284/*284:xpc10:284*/;
           A_SINT[19'h6_1fe8+9'h1b8] <= -32'd3;
           end 
          
      9'd284/*284:US*/:  begin 
           xpc10 <= 9'd285/*285:xpc10:285*/;
           A_SINT[19'h6_1fe8+9'h1bc] <= 32'd0;
           end 
          
      9'd285/*285:US*/:  begin 
           xpc10 <= 9'd286/*286:xpc10:286*/;
           A_SINT[19'h6_1fe8+9'h1c0] <= -32'd1;
           end 
          
      9'd286/*286:US*/:  begin 
           xpc10 <= 9'd287/*287:xpc10:287*/;
           A_SINT[19'h6_1fe8+9'h1c4] <= -32'd1;
           end 
          
      9'd287/*287:US*/:  begin 
           xpc10 <= 9'd288/*288:xpc10:288*/;
           A_SINT[19'h6_1fe8+9'h1c8] <= -32'd3;
           end 
          
      9'd288/*288:US*/:  begin 
           xpc10 <= 9'd289/*289:xpc10:289*/;
           A_SINT[19'h6_1fe8+9'h1cc] <= 32'd1;
           end 
          
      9'd289/*289:US*/:  begin 
           xpc10 <= 9'd290/*290:xpc10:290*/;
           A_SINT[19'h6_1fe8+9'h1d0] <= 32'd0;
           end 
          
      9'd290/*290:US*/:  begin 
           xpc10 <= 9'd291/*291:xpc10:291*/;
           A_SINT[19'h6_1fe8+9'h1d4] <= -32'd1;
           end 
          
      9'd291/*291:US*/:  begin 
           xpc10 <= 9'd292/*292:xpc10:292*/;
           A_SINT[19'h6_1fe8+9'h1d8] <= -32'd7;
           end 
          
      9'd292/*292:US*/:  begin 
           xpc10 <= 9'd293/*293:xpc10:293*/;
           A_SINT[19'h6_1fe8+9'h1dc] <= -32'd5;
           end 
          
      9'd293/*293:US*/:  begin 
           xpc10 <= 9'd294/*294:xpc10:294*/;
           A_SINT[19'h6_1fe8+9'h1e0] <= -32'd1;
           end 
          
      9'd294/*294:US*/:  begin 
           xpc10 <= 9'd295/*295:xpc10:295*/;
           A_SINT[19'h6_1fe8+9'h1e4] <= -32'd3;
           end 
          
      9'd295/*295:US*/:  begin 
           xpc10 <= 9'd296/*296:xpc10:296*/;
           A_SINT[19'h6_1fe8+9'h1e8] <= 32'd1;
           end 
          
      9'd296/*296:US*/:  begin 
           xpc10 <= 9'd297/*297:xpc10:297*/;
           A_SINT[19'h6_1fe8+9'h1ec] <= 32'd1;
           end 
          
      9'd297/*297:US*/:  begin 
           xpc10 <= 9'd298/*298:xpc10:298*/;
           A_SINT[19'h6_1fe8+9'h1f0] <= -32'd2;
           end 
          
      9'd298/*298:US*/:  begin 
           xpc10 <= 9'd299/*299:xpc10:299*/;
           A_SINT[19'h6_1fe8+9'h1f4] <= -32'd2;
           end 
          
      9'd299/*299:US*/:  begin 
           xpc10 <= 9'd300/*300:xpc10:300*/;
           A_SINT[19'h6_1fe8+9'h1f8] <= 32'd6;
           end 
          
      9'd300/*300:US*/:  begin 
           xpc10 <= 9'd301/*301:xpc10:301*/;
           A_SINT[19'h6_1fe8+9'h1fc] <= -32'd2;
           end 
          
      9'd301/*301:US*/:  begin 
           xpc10 <= 9'd302/*302:xpc10:302*/;
           A_SINT[19'h6_1fe8+10'h200] <= 32'd0;
           end 
          
      9'd302/*302:US*/:  begin 
           xpc10 <= 9'd303/*303:xpc10:303*/;
           A_SINT[19'h6_1fe8+10'h204] <= -32'd2;
           end 
          
      9'd303/*303:US*/:  begin 
           xpc10 <= 9'd304/*304:xpc10:304*/;
           A_SINT[19'h6_1fe8+10'h208] <= -32'd2;
           end 
          
      9'd304/*304:US*/:  begin 
           xpc10 <= 9'd305/*305:xpc10:305*/;
           A_SINT[19'h6_1fe8+10'h20c] <= 32'd2;
           end 
          
      9'd305/*305:US*/:  begin 
           xpc10 <= 9'd306/*306:xpc10:306*/;
           A_SINT[19'h6_1fe8+10'h210] <= 32'd0;
           end 
          
      9'd306/*306:US*/:  begin 
           xpc10 <= 9'd307/*307:xpc10:307*/;
           A_SINT[19'h6_1fe8+10'h214] <= 32'd3;
           end 
          
      9'd307/*307:US*/:  begin 
           xpc10 <= 9'd308/*308:xpc10:308*/;
           A_SINT[19'h6_1fe8+10'h218] <= 32'd2;
           end 
          
      9'd308/*308:US*/:  begin 
           xpc10 <= 9'd309/*309:xpc10:309*/;
           A_SINT[19'h6_1fe8+10'h21c] <= -32'd1;
           end 
          
      9'd309/*309:US*/:  begin 
           xpc10 <= 9'd310/*310:xpc10:310*/;
           A_SINT[19'h6_1fe8+10'h220] <= -32'd1;
           end 
          
      9'd310/*310:US*/:  begin 
           xpc10 <= 9'd311/*311:xpc10:311*/;
           A_SINT[19'h6_1fe8+10'h224] <= -32'd2;
           end 
          
      9'd311/*311:US*/:  begin 
           xpc10 <= 9'd312/*312:xpc10:312*/;
           A_SINT[19'h6_1fe8+10'h228] <= -32'd3;
           end 
          
      9'd312/*312:US*/:  begin 
           xpc10 <= 9'd313/*313:xpc10:313*/;
           A_SINT[19'h6_1fe8+10'h22c] <= 32'd0;
           end 
          
      9'd313/*313:US*/:  begin 
           xpc10 <= 9'd314/*314:xpc10:314*/;
           A_SINT[19'h6_1fe8+10'h230] <= -32'd1;
           end 
          
      9'd314/*314:US*/:  begin 
           xpc10 <= 9'd315/*315:xpc10:315*/;
           A_SINT[19'h6_1fe8+10'h234] <= -32'd2;
           end 
          
      9'd315/*315:US*/:  begin 
           xpc10 <= 9'd316/*316:xpc10:316*/;
           A_SINT[19'h6_1fe8+10'h238] <= -32'd2;
           end 
          
      9'd316/*316:US*/:  begin 
           xpc10 <= 9'd317/*317:xpc10:317*/;
           A_SINT[19'h6_1fe8+10'h23c] <= -32'd2;
           end 
          
      9'd317/*317:US*/:  begin 
           xpc10 <= 9'd318/*318:xpc10:318*/;
           A_SINT[19'h6_1fe8+10'h240] <= 32'd1;
           end 
          
      9'd318/*318:US*/:  begin 
           xpc10 <= 9'd319/*319:xpc10:319*/;
           A_SINT[19'h6_1fe8+10'h244] <= -32'd3;
           end 
          
      9'd319/*319:US*/:  begin 
           xpc10 <= 9'd320/*320:xpc10:320*/;
           A_SINT[19'h6_1fe8+10'h248] <= -32'd2;
           end 
          
      9'd320/*320:US*/:  begin 
           xpc10 <= 9'd321/*321:xpc10:321*/;
           A_SINT[19'h6_1fe8+10'h24c] <= 32'd5;
           end 
          
      9'd321/*321:US*/:  begin 
           xpc10 <= 9'd322/*322:xpc10:322*/;
           A_SINT[19'h6_1fe8+10'h250] <= -32'd2;
           end 
          
      9'd322/*322:US*/:  begin 
           xpc10 <= 9'd323/*323:xpc10:323*/;
           A_SINT[19'h6_1fe8+10'h254] <= 32'd2;
           end 
          
      9'd323/*323:US*/:  begin 
           xpc10 <= 9'd324/*324:xpc10:324*/;
           A_SINT[19'h6_1fe8+10'h258] <= 32'd2;
           end 
          
      9'd324/*324:US*/:  begin 
           xpc10 <= 9'd325/*325:xpc10:325*/;
           A_SINT[19'h6_1fe8+10'h25c] <= -32'd2;
           end 
          
      9'd325/*325:US*/:  begin 
           xpc10 <= 9'd326/*326:xpc10:326*/;
           A_SINT[19'h6_1fe8+10'h260] <= -32'd2;
           end 
          
      9'd326/*326:US*/:  begin 
           xpc10 <= 9'd327/*327:xpc10:327*/;
           A_SINT[19'h6_1fe8+10'h264] <= -32'd2;
           end 
          
      9'd327/*327:US*/:  begin 
           xpc10 <= 9'd328/*328:xpc10:328*/;
           A_SINT[19'h6_1fe8+10'h268] <= -32'd2;
           end 
          
      9'd328/*328:US*/:  begin 
           xpc10 <= 9'd329/*329:xpc10:329*/;
           A_SINT[19'h6_1fe8+10'h26c] <= -32'd1;
           end 
          
      9'd329/*329:US*/:  begin 
           xpc10 <= 9'd330/*330:xpc10:330*/;
           A_SINT[19'h6_1fe8+10'h270] <= 32'd0;
           end 
          
      9'd330/*330:US*/:  begin 
           xpc10 <= 9'd331/*331:xpc10:331*/;
           A_SINT[19'h6_1fe8+10'h274] <= 32'd4;
           end 
          
      9'd331/*331:US*/:  begin 
           xpc10 <= 9'd332/*332:xpc10:332*/;
           A_SINT[19'h6_1fe8+10'h278] <= -32'd5;
           end 
          
      9'd332/*332:US*/:  begin 
           xpc10 <= 9'd333/*333:xpc10:333*/;
           A_SINT[19'h6_1fe8+10'h27c] <= -32'd1;
           end 
          
      9'd333/*333:US*/:  begin 
           xpc10 <= 9'd334/*334:xpc10:334*/;
           A_SINT[19'h6_1fe8+10'h280] <= -32'd1;
           end 
          
      9'd334/*334:US*/:  begin 
           xpc10 <= 9'd335/*335:xpc10:335*/;
           A_SINT[19'h6_1fe8+10'h284] <= -32'd5;
           end 
          
      9'd335/*335:US*/:  begin 
           xpc10 <= 9'd336/*336:xpc10:336*/;
           A_SINT[19'h6_1fe8+10'h288] <= 32'd0;
           end 
          
      9'd336/*336:US*/:  begin 
           xpc10 <= 9'd337/*337:xpc10:337*/;
           A_SINT[19'h6_1fe8+10'h28c] <= 32'd0;
           end 
          
      9'd337/*337:US*/:  begin 
           xpc10 <= 9'd338/*338:xpc10:338*/;
           A_SINT[19'h6_1fe8+10'h290] <= -32'd5;
           end 
          
      9'd338/*338:US*/:  begin 
           xpc10 <= 9'd339/*339:xpc10:339*/;
           A_SINT[19'h6_1fe8+10'h294] <= -32'd2;
           end 
          
      9'd339/*339:US*/:  begin 
           xpc10 <= 9'd340/*340:xpc10:340*/;
           A_SINT[19'h6_1fe8+10'h298] <= 32'd0;
           end 
          
      9'd340/*340:US*/:  begin 
           xpc10 <= 9'd341/*341:xpc10:341*/;
           A_SINT[19'h6_1fe8+10'h29c] <= -32'd2;
           end 
          
      9'd341/*341:US*/:  begin 
           xpc10 <= 9'd342/*342:xpc10:342*/;
           A_SINT[19'h6_1fe8+10'h2a0] <= 32'd5;
           end 
          
      9'd342/*342:US*/:  begin 
           xpc10 <= 9'd343/*343:xpc10:343*/;
           A_SINT[19'h6_1fe8+10'h2a4] <= -32'd3;
           end 
          
      9'd343/*343:US*/:  begin 
           xpc10 <= 9'd344/*344:xpc10:344*/;
           A_SINT[19'h6_1fe8+10'h2a8] <= 32'd0;
           end 
          
      9'd344/*344:US*/:  begin 
           xpc10 <= 9'd345/*345:xpc10:345*/;
           A_SINT[19'h6_1fe8+10'h2ac] <= 32'd1;
           end 
          
      9'd345/*345:US*/:  begin 
           xpc10 <= 9'd346/*346:xpc10:346*/;
           A_SINT[19'h6_1fe8+10'h2b0] <= -32'd1;
           end 
          
      9'd346/*346:US*/:  begin 
           xpc10 <= 9'd347/*347:xpc10:347*/;
           A_SINT[19'h6_1fe8+10'h2b4] <= 32'd1;
           end 
          
      9'd347/*347:US*/:  begin 
           xpc10 <= 9'd348/*348:xpc10:348*/;
           A_SINT[19'h6_1fe8+10'h2b8] <= 32'd3;
           end 
          
      9'd348/*348:US*/:  begin 
           xpc10 <= 9'd349/*349:xpc10:349*/;
           A_SINT[19'h6_1fe8+10'h2bc] <= 32'd0;
           end 
          
      9'd349/*349:US*/:  begin 
           xpc10 <= 9'd350/*350:xpc10:350*/;
           A_SINT[19'h6_1fe8+10'h2c0] <= 32'd0;
           end 
          
      9'd350/*350:US*/:  begin 
           xpc10 <= 9'd351/*351:xpc10:351*/;
           A_SINT[19'h6_1fe8+10'h2c4] <= -32'd2;
           end 
          
      9'd351/*351:US*/:  begin 
           xpc10 <= 9'd352/*352:xpc10:352*/;
           A_SINT[19'h6_1fe8+10'h2c8] <= -32'd3;
           end 
          
      9'd352/*352:US*/:  begin 
           xpc10 <= 9'd353/*353:xpc10:353*/;
           A_SINT[19'h6_1fe8+10'h2cc] <= -32'd4;
           end 
          
      9'd353/*353:US*/:  begin 
           xpc10 <= 9'd354/*354:xpc10:354*/;
           A_SINT[19'h6_1fe8+10'h2d0] <= -32'd2;
           end 
          
      9'd354/*354:US*/:  begin 
           xpc10 <= 9'd355/*355:xpc10:355*/;
           A_SINT[19'h6_1fe8+10'h2d4] <= -32'd6;
           end 
          
      9'd355/*355:US*/:  begin 
           xpc10 <= 9'd356/*356:xpc10:356*/;
           A_SINT[19'h6_1fe8+10'h2d8] <= -32'd4;
           end 
          
      9'd356/*356:US*/:  begin 
           xpc10 <= 9'd357/*357:xpc10:357*/;
           A_SINT[19'h6_1fe8+10'h2dc] <= -32'd3;
           end 
          
      9'd357/*357:US*/:  begin 
           xpc10 <= 9'd358/*358:xpc10:358*/;
           A_SINT[19'h6_1fe8+10'h2e0] <= 32'd2;
           end 
          
      9'd358/*358:US*/:  begin 
           xpc10 <= 9'd359/*359:xpc10:359*/;
           A_SINT[19'h6_1fe8+10'h2e4] <= -32'd4;
           end 
          
      9'd359/*359:US*/:  begin 
           xpc10 <= 9'd360/*360:xpc10:360*/;
           A_SINT[19'h6_1fe8+10'h2e8] <= -32'd2;
           end 
          
      9'd360/*360:US*/:  begin 
           xpc10 <= 9'd361/*361:xpc10:361*/;
           A_SINT[19'h6_1fe8+10'h2ec] <= 32'd2;
           end 
          
      9'd361/*361:US*/:  begin 
           xpc10 <= 9'd362/*362:xpc10:362*/;
           A_SINT[19'h6_1fe8+10'h2f0] <= -32'd3;
           end 
          
      9'd362/*362:US*/:  begin 
           xpc10 <= 9'd363/*363:xpc10:363*/;
           A_SINT[19'h6_1fe8+10'h2f4] <= 32'd6;
           end 
          
      9'd363/*363:US*/:  begin 
           xpc10 <= 9'd364/*364:xpc10:364*/;
           A_SINT[19'h6_1fe8+10'h2f8] <= 32'd4;
           end 
          
      9'd364/*364:US*/:  begin 
           xpc10 <= 9'd365/*365:xpc10:365*/;
           A_SINT[19'h6_1fe8+10'h2fc] <= -32'd3;
           end 
          
      9'd365/*365:US*/:  begin 
           xpc10 <= 9'd366/*366:xpc10:366*/;
           A_SINT[19'h6_1fe8+10'h300] <= -32'd3;
           end 
          
      9'd366/*366:US*/:  begin 
           xpc10 <= 9'd367/*367:xpc10:367*/;
           A_SINT[19'h6_1fe8+10'h304] <= -32'd2;
           end 
          
      9'd367/*367:US*/:  begin 
           xpc10 <= 9'd368/*368:xpc10:368*/;
           A_SINT[19'h6_1fe8+10'h308] <= -32'd3;
           end 
          
      9'd368/*368:US*/:  begin 
           xpc10 <= 9'd369/*369:xpc10:369*/;
           A_SINT[19'h6_1fe8+10'h30c] <= -32'd3;
           end 
          
      9'd369/*369:US*/:  begin 
           xpc10 <= 9'd370/*370:xpc10:370*/;
           A_SINT[19'h6_1fe8+10'h310] <= -32'd2;
           end 
          
      9'd370/*370:US*/:  begin 
           xpc10 <= 9'd371/*371:xpc10:371*/;
           A_SINT[19'h6_1fe8+10'h314] <= 32'd2;
           end 
          
      9'd371/*371:US*/:  begin 
           xpc10 <= 9'd372/*372:xpc10:372*/;
           A_SINT[19'h6_1fe8+10'h318] <= -32'd2;
           end 
          
      9'd372/*372:US*/:  begin 
           xpc10 <= 9'd373/*373:xpc10:373*/;
           A_SINT[19'h6_1fe8+10'h31c] <= -32'd1;
           end 
          
      9'd373/*373:US*/:  begin 
           xpc10 <= 9'd374/*374:xpc10:374*/;
           A_SINT[19'h6_1fe8+10'h320] <= -32'd1;
           end 
          
      9'd374/*374:US*/:  begin 
           xpc10 <= 9'd375/*375:xpc10:375*/;
           A_SINT[19'h6_1fe8+10'h324] <= -32'd5;
           end 
          
      9'd375/*375:US*/:  begin 
           xpc10 <= 9'd376/*376:xpc10:376*/;
           A_SINT[19'h6_1fe8+10'h328] <= -32'd3;
           end 
          
      9'd376/*376:US*/:  begin 
           xpc10 <= 9'd377/*377:xpc10:377*/;
           A_SINT[19'h6_1fe8+10'h32c] <= -32'd2;
           end 
          
      9'd377/*377:US*/:  begin 
           xpc10 <= 9'd378/*378:xpc10:378*/;
           A_SINT[19'h6_1fe8+10'h330] <= 32'd0;
           end 
          
      9'd378/*378:US*/:  begin 
           xpc10 <= 9'd379/*379:xpc10:379*/;
           A_SINT[19'h6_1fe8+10'h334] <= -32'd3;
           end 
          
      9'd379/*379:US*/:  begin 
           xpc10 <= 9'd380/*380:xpc10:380*/;
           A_SINT[19'h6_1fe8+10'h338] <= -32'd2;
           end 
          
      9'd380/*380:US*/:  begin 
           xpc10 <= 9'd381/*381:xpc10:381*/;
           A_SINT[19'h6_1fe8+10'h33c] <= 32'd2;
           end 
          
      9'd381/*381:US*/:  begin 
           xpc10 <= 9'd382/*382:xpc10:382*/;
           A_SINT[19'h6_1fe8+10'h340] <= 32'd0;
           end 
          
      9'd382/*382:US*/:  begin 
           xpc10 <= 9'd383/*383:xpc10:383*/;
           A_SINT[19'h6_1fe8+10'h344] <= 32'd4;
           end 
          
      9'd383/*383:US*/:  begin 
           xpc10 <= 9'd384/*384:xpc10:384*/;
           A_SINT[19'h6_1fe8+10'h348] <= 32'd6;
           end 
          
      9'd384/*384:US*/:  begin 
           xpc10 <= 9'd385/*385:xpc10:385*/;
           A_SINT[19'h6_1fe8+10'h34c] <= -32'd2;
           end 
          
      9'd385/*385:US*/:  begin 
           xpc10 <= 9'd386/*386:xpc10:386*/;
           A_SINT[19'h6_1fe8+10'h350] <= -32'd2;
           end 
          
      9'd386/*386:US*/:  begin 
           xpc10 <= 9'd387/*387:xpc10:387*/;
           A_SINT[19'h6_1fe8+10'h354] <= -32'd1;
           end 
          
      9'd387/*387:US*/:  begin 
           xpc10 <= 9'd388/*388:xpc10:388*/;
           A_SINT[19'h6_1fe8+10'h358] <= 32'd0;
           end 
          
      9'd388/*388:US*/:  begin 
           xpc10 <= 9'd389/*389:xpc10:389*/;
           A_SINT[19'h6_1fe8+10'h35c] <= -32'd2;
           end 
          
      9'd389/*389:US*/:  begin 
           xpc10 <= 9'd390/*390:xpc10:390*/;
           A_SINT[19'h6_1fe8+10'h360] <= -32'd1;
           end 
          
      9'd390/*390:US*/:  begin 
           xpc10 <= 9'd391/*391:xpc10:391*/;
           A_SINT[19'h6_1fe8+10'h364] <= 32'd2;
           end 
          
      9'd391/*391:US*/:  begin 
           xpc10 <= 9'd392/*392:xpc10:392*/;
           A_SINT[19'h6_1fe8+10'h368] <= -32'd4;
           end 
          
      9'd392/*392:US*/:  begin 
           xpc10 <= 9'd393/*393:xpc10:393*/;
           A_SINT[19'h6_1fe8+10'h36c] <= -32'd2;
           end 
          
      9'd393/*393:US*/:  begin 
           xpc10 <= 9'd394/*394:xpc10:394*/;
           A_SINT[19'h6_1fe8+10'h370] <= 32'd0;
           end 
          
      9'd394/*394:US*/:  begin 
           xpc10 <= 9'd395/*395:xpc10:395*/;
           A_SINT[19'h6_1fe8+10'h374] <= -32'd4;
           end 
          
      9'd395/*395:US*/:  begin 
           xpc10 <= 9'd396/*396:xpc10:396*/;
           A_SINT[19'h6_1fe8+10'h378] <= 32'd2;
           end 
          
      9'd396/*396:US*/:  begin 
           xpc10 <= 9'd397/*397:xpc10:397*/;
           A_SINT[19'h6_1fe8+10'h37c] <= 32'd1;
           end 
          
      9'd397/*397:US*/:  begin 
           xpc10 <= 9'd398/*398:xpc10:398*/;
           A_SINT[19'h6_1fe8+10'h380] <= -32'd4;
           end 
          
      9'd398/*398:US*/:  begin 
           xpc10 <= 9'd399/*399:xpc10:399*/;
           A_SINT[19'h6_1fe8+10'h384] <= 32'd0;
           end 
          
      9'd399/*399:US*/:  begin 
           xpc10 <= 9'd400/*400:xpc10:400*/;
           A_SINT[19'h6_1fe8+10'h388] <= 32'd2;
           end 
          
      9'd400/*400:US*/:  begin 
           xpc10 <= 9'd401/*401:xpc10:401*/;
           A_SINT[19'h6_1fe8+10'h38c] <= -32'd2;
           end 
          
      9'd401/*401:US*/:  begin 
           xpc10 <= 9'd402/*402:xpc10:402*/;
           A_SINT[19'h6_1fe8+10'h390] <= 32'd1;
           end 
          
      9'd402/*402:US*/:  begin 
           xpc10 <= 9'd403/*403:xpc10:403*/;
           A_SINT[19'h6_1fe8+10'h394] <= -32'd3;
           end 
          
      9'd403/*403:US*/:  begin 
           xpc10 <= 9'd404/*404:xpc10:404*/;
           A_SINT[19'h6_1fe8+10'h398] <= -32'd2;
           end 
          
      9'd404/*404:US*/:  begin 
           xpc10 <= 9'd405/*405:xpc10:405*/;
           A_SINT[19'h6_1fe8+10'h39c] <= 32'd2;
           end 
          
      9'd405/*405:US*/:  begin 
           xpc10 <= 9'd406/*406:xpc10:406*/;
           A_SINT[19'h6_1fe8+10'h3a0] <= -32'd1;
           end 
          
      9'd406/*406:US*/:  begin 
           xpc10 <= 9'd407/*407:xpc10:407*/;
           A_SINT[19'h6_1fe8+10'h3a4] <= 32'd1;
           end 
          
      9'd407/*407:US*/:  begin 
           xpc10 <= 9'd408/*408:xpc10:408*/;
           A_SINT[19'h6_1fe8+10'h3a8] <= 32'd0;
           end 
          
      9'd408/*408:US*/:  begin 
           xpc10 <= 9'd409/*409:xpc10:409*/;
           A_SINT[19'h6_1fe8+10'h3ac] <= 32'd1;
           end 
          
      9'd409/*409:US*/:  begin 
           xpc10 <= 9'd410/*410:xpc10:410*/;
           A_SINT[19'h6_1fe8+10'h3b0] <= 32'd0;
           end 
          
      9'd410/*410:US*/:  begin 
           xpc10 <= 9'd411/*411:xpc10:411*/;
           A_SINT[19'h6_1fe8+10'h3b4] <= -32'd2;
           end 
          
      9'd411/*411:US*/:  begin 
           xpc10 <= 9'd412/*412:xpc10:412*/;
           A_SINT[19'h6_1fe8+10'h3b8] <= -32'd4;
           end 
          
      9'd412/*412:US*/:  begin 
           xpc10 <= 9'd413/*413:xpc10:413*/;
           A_SINT[19'h6_1fe8+10'h3bc] <= -32'd2;
           end 
          
      9'd413/*413:US*/:  begin 
           xpc10 <= 9'd414/*414:xpc10:414*/;
           A_SINT[19'h6_1fe8+10'h3c0] <= 32'd1;
           end 
          
      9'd414/*414:US*/:  begin 
           xpc10 <= 9'd415/*415:xpc10:415*/;
           A_SINT[19'h6_1fe8+10'h3c4] <= -32'd3;
           end 
          
      9'd415/*415:US*/:  begin 
           xpc10 <= 9'd416/*416:xpc10:416*/;
           A_SINT[19'h6_1fe8+10'h3c8] <= -32'd1;
           end 
          
      9'd416/*416:US*/:  begin 
           xpc10 <= 9'd417/*417:xpc10:417*/;
           A_SINT[19'h6_1fe8+10'h3cc] <= -32'd1;
           end 
          
      9'd417/*417:US*/:  begin 
           xpc10 <= 9'd418/*418:xpc10:418*/;
           A_SINT[19'h6_1fe8+10'h3d0] <= -32'd5;
           end 
          
      9'd418/*418:US*/:  begin 
           xpc10 <= 9'd419/*419:xpc10:419*/;
           A_SINT[19'h6_1fe8+10'h3d4] <= -32'd1;
           end 
          
      9'd419/*419:US*/:  begin 
           xpc10 <= 9'd420/*420:xpc10:420*/;
           A_SINT[19'h6_1fe8+10'h3d8] <= 32'd0;
           end 
          
      9'd420/*420:US*/:  begin 
           xpc10 <= 9'd421/*421:xpc10:421*/;
           A_SINT[19'h6_1fe8+10'h3dc] <= -32'd2;
           end 
          
      9'd421/*421:US*/:  begin 
           xpc10 <= 9'd422/*422:xpc10:422*/;
           A_SINT[19'h6_1fe8+10'h3e0] <= -32'd1;
           end 
          
      9'd422/*422:US*/:  begin 
           xpc10 <= 9'd423/*423:xpc10:423*/;
           A_SINT[19'h6_1fe8+10'h3e4] <= -32'd3;
           end 
          
      9'd423/*423:US*/:  begin 
           xpc10 <= 9'd424/*424:xpc10:424*/;
           A_SINT[19'h6_1fe8+10'h3e8] <= -32'd2;
           end 
          
      9'd424/*424:US*/:  begin 
           xpc10 <= 9'd425/*425:xpc10:425*/;
           A_SINT[19'h6_1fe8+10'h3ec] <= -32'd1;
           end 
          
      9'd425/*425:US*/:  begin 
           xpc10 <= 9'd426/*426:xpc10:426*/;
           A_SINT[19'h6_1fe8+10'h3f0] <= 32'd6;
           end 
          
      9'd426/*426:US*/:  begin 
           xpc10 <= 9'd427/*427:xpc10:427*/;
           A_SINT[19'h6_1fe8+10'h3f4] <= 32'd0;
           end 
          
      9'd427/*427:US*/:  begin 
           xpc10 <= 9'd428/*428:xpc10:428*/;
           A_SINT[19'h6_1fe8+10'h3f8] <= 32'd0;
           end 
          
      9'd428/*428:US*/:  begin 
           xpc10 <= 9'd429/*429:xpc10:429*/;
           A_SINT[19'h6_1fe8+10'h3fc] <= 32'd1;
           end 
          
      9'd429/*429:US*/:  begin 
           xpc10 <= 9'd430/*430:xpc10:430*/;
           A_SINT[19'h6_1fe8+11'h400] <= 32'd0;
           end 
          
      9'd430/*430:US*/:  begin 
           xpc10 <= 9'd431/*431:xpc10:431*/;
           A_SINT[19'h6_1fe8+11'h404] <= -32'd1;
           end 
          
      9'd431/*431:US*/:  begin 
           xpc10 <= 9'd432/*432:xpc10:432*/;
           A_SINT[19'h6_1fe8+11'h408] <= -32'd6;
           end 
          
      9'd432/*432:US*/:  begin 
           xpc10 <= 9'd433/*433:xpc10:433*/;
           A_SINT[19'h6_1fe8+11'h40c] <= -32'd5;
           end 
          
      9'd433/*433:US*/:  begin 
           xpc10 <= 9'd434/*434:xpc10:434*/;
           A_SINT[19'h6_1fe8+11'h410] <= 32'd0;
           end 
          
      9'd434/*434:US*/:  begin 
           xpc10 <= 9'd435/*435:xpc10:435*/;
           A_SINT[19'h6_1fe8+11'h414] <= -32'd5;
           end 
          
      9'd435/*435:US*/:  begin 
           xpc10 <= 9'd436/*436:xpc10:436*/;
           A_SINT[19'h6_1fe8+11'h418] <= 32'd2;
           end 
          
      9'd436/*436:US*/:  begin 
           xpc10 <= 9'd437/*437:xpc10:437*/;
           A_SINT[19'h6_1fe8+11'h41c] <= 32'd2;
           end 
          
      9'd437/*437:US*/:  begin 
           xpc10 <= 9'd438/*438:xpc10:438*/;
           A_SINT[19'h6_1fe8+11'h420] <= -32'd5;
           end 
          
      9'd438/*438:US*/:  begin 
           xpc10 <= 9'd439/*439:xpc10:439*/;
           A_SINT[19'h6_1fe8+11'h424] <= -32'd1;
           end 
          
      9'd439/*439:US*/:  begin 
           xpc10 <= 9'd440/*440:xpc10:440*/;
           A_SINT[19'h6_1fe8+11'h428] <= 32'd3;
           end 
          
      9'd440/*440:US*/:  begin 
           xpc10 <= 9'd441/*441:xpc10:441*/;
           A_SINT[19'h6_1fe8+11'h42c] <= -32'd2;
           end 
          
      9'd441/*441:US*/:  begin 
           xpc10 <= 9'd442/*442:xpc10:442*/;
           A_SINT[19'h6_1fe8+11'h430] <= 32'd1;
           end 
          
      9'd442/*442:US*/:  begin 
           xpc10 <= 9'd443/*443:xpc10:443*/;
           A_SINT[19'h6_1fe8+11'h434] <= -32'd2;
           end 
          
      9'd443/*443:US*/:  begin 
           xpc10 <= 9'd444/*444:xpc10:444*/;
           A_SINT[19'h6_1fe8+11'h438] <= -32'd1;
           end 
          
      9'd444/*444:US*/:  begin 
           xpc10 <= 9'd445/*445:xpc10:445*/;
           A_SINT[19'h6_1fe8+11'h43c] <= 32'd1;
           end 
          
      9'd445/*445:US*/:  begin 
           xpc10 <= 9'd446/*446:xpc10:446*/;
           A_SINT[19'h6_1fe8+11'h440] <= 32'd0;
           end 
          
      9'd446/*446:US*/:  begin 
           xpc10 <= 9'd447/*447:xpc10:447*/;
           A_SINT[19'h6_1fe8+11'h444] <= 32'd4;
           end 
          
      9'd447/*447:US*/:  begin 
           xpc10 <= 9'd448/*448:xpc10:448*/;
           A_SINT[19'h6_1fe8+11'h448] <= 32'd1;
           end 
          
      9'd448/*448:US*/:  begin 
           xpc10 <= 9'd449/*449:xpc10:449*/;
           A_SINT[19'h6_1fe8+11'h44c] <= -32'd1;
           end 
          
      9'd449/*449:US*/:  begin 
           xpc10 <= 9'd450/*450:xpc10:450*/;
           A_SINT[19'h6_1fe8+11'h450] <= -32'd1;
           end 
          
      9'd450/*450:US*/:  begin 
           xpc10 <= 9'd451/*451:xpc10:451*/;
           A_SINT[19'h6_1fe8+11'h454] <= -32'd2;
           end 
          
      9'd451/*451:US*/:  begin 
           xpc10 <= 9'd452/*452:xpc10:452*/;
           A_SINT[19'h6_1fe8+11'h458] <= -32'd5;
           end 
          
      9'd452/*452:US*/:  begin 
           xpc10 <= 9'd453/*453:xpc10:453*/;
           A_SINT[19'h6_1fe8+11'h45c] <= -32'd4;
           end 
          
      9'd453/*453:US*/:  begin 
           xpc10 <= 9'd454/*454:xpc10:454*/;
           A_SINT[19'h6_1fe8+11'h460] <= -32'd2;
           end 
          
      9'd454/*454:US*/:  begin 
           xpc10 <= 9'd455/*455:xpc10:455*/;
           A_SINT[19'h6_1fe8+11'h464] <= -32'd4;
           end 
          
      9'd455/*455:US*/:  begin 
           xpc10 <= 9'd456/*456:xpc10:456*/;
           A_SINT[19'h6_1fe8+11'h468] <= -32'd1;
           end 
          
      9'd456/*456:US*/:  begin 
           xpc10 <= 9'd457/*457:xpc10:457*/;
           A_SINT[19'h6_1fe8+11'h46c] <= -32'd1;
           end 
          
      9'd457/*457:US*/:  begin 
           xpc10 <= 9'd458/*458:xpc10:458*/;
           A_SINT[19'h6_1fe8+11'h470] <= -32'd4;
           end 
          
      9'd458/*458:US*/:  begin 
           xpc10 <= 9'd459/*459:xpc10:459*/;
           A_SINT[19'h6_1fe8+11'h474] <= -32'd3;
           end 
          
      9'd459/*459:US*/:  begin 
           xpc10 <= 9'd460/*460:xpc10:460*/;
           A_SINT[19'h6_1fe8+11'h478] <= 32'd2;
           end 
          
      9'd460/*460:US*/:  begin 
           xpc10 <= 9'd461/*461:xpc10:461*/;
           A_SINT[19'h6_1fe8+11'h47c] <= -32'd2;
           end 
          
      9'd461/*461:US*/:  begin 
           xpc10 <= 9'd462/*462:xpc10:462*/;
           A_SINT[19'h6_1fe8+11'h480] <= 32'd3;
           end 
          
      9'd462/*462:US*/:  begin 
           xpc10 <= 9'd463/*463:xpc10:463*/;
           A_SINT[19'h6_1fe8+11'h484] <= -32'd3;
           end 
          
      9'd463/*463:US*/:  begin 
           xpc10 <= 9'd464/*464:xpc10:464*/;
           A_SINT[19'h6_1fe8+11'h488] <= 32'd0;
           end 
          
      9'd464/*464:US*/:  begin 
           xpc10 <= 9'd465/*465:xpc10:465*/;
           A_SINT[19'h6_1fe8+11'h48c] <= 32'd0;
           end 
          
      9'd465/*465:US*/:  begin 
           xpc10 <= 9'd466/*466:xpc10:466*/;
           A_SINT[19'h6_1fe8+11'h490] <= 32'd0;
           end 
          
      9'd466/*466:US*/:  begin 
           xpc10 <= 9'd467/*467:xpc10:467*/;
           A_SINT[19'h6_1fe8+11'h494] <= 32'd1;
           end 
          
      9'd467/*467:US*/:  begin 
           xpc10 <= 9'd468/*468:xpc10:468*/;
           A_SINT[19'h6_1fe8+11'h498] <= 32'd6;
           end 
          
      9'd468/*468:US*/:  begin 
           xpc10 <= 9'd469/*469:xpc10:469*/;
           A_SINT[19'h6_1fe8+11'h49c] <= 32'd0;
           end 
          
      9'd469/*469:US*/:  begin 
           xpc10 <= 9'd470/*470:xpc10:470*/;
           A_SINT[19'h6_1fe8+11'h4a0] <= -32'd1;
           end 
          
      9'd470/*470:US*/:  begin 
           xpc10 <= 9'd471/*471:xpc10:471*/;
           A_SINT[19'h6_1fe8+11'h4a4] <= -32'd2;
           end 
          
      9'd471/*471:US*/:  begin 
           xpc10 <= 9'd472/*472:xpc10:472*/;
           A_SINT[19'h6_1fe8+11'h4a8] <= 32'd2;
           end 
          
      9'd472/*472:US*/:  begin 
           xpc10 <= 9'd473/*473:xpc10:473*/;
           A_SINT[19'h6_1fe8+11'h4ac] <= -32'd4;
           end 
          
      9'd473/*473:US*/:  begin 
           xpc10 <= 9'd474/*474:xpc10:474*/;
           A_SINT[19'h6_1fe8+11'h4b0] <= 32'd1;
           end 
          
      9'd474/*474:US*/:  begin 
           xpc10 <= 9'd475/*475:xpc10:475*/;
           A_SINT[19'h6_1fe8+11'h4b4] <= 32'd0;
           end 
          
      9'd475/*475:US*/:  begin 
           xpc10 <= 9'd476/*476:xpc10:476*/;
           A_SINT[19'h6_1fe8+11'h4b8] <= 32'd0;
           end 
          
      9'd476/*476:US*/:  begin 
           xpc10 <= 9'd477/*477:xpc10:477*/;
           A_SINT[19'h6_1fe8+11'h4bc] <= 32'd0;
           end 
          
      9'd477/*477:US*/:  begin 
           xpc10 <= 9'd478/*478:xpc10:478*/;
           A_SINT[19'h6_1fe8+11'h4c0] <= -32'd3;
           end 
          
      9'd478/*478:US*/:  begin 
           xpc10 <= 9'd479/*479:xpc10:479*/;
           A_SINT[19'h6_1fe8+11'h4c4] <= 32'd1;
           end 
          
      9'd479/*479:US*/:  begin 
           xpc10 <= 9'd480/*480:xpc10:480*/;
           A_SINT[19'h6_1fe8+11'h4c8] <= -32'd1;
           end 
          
      9'd480/*480:US*/:  begin 
           xpc10 <= 9'd481/*481:xpc10:481*/;
           A_SINT[19'h6_1fe8+11'h4cc] <= -32'd1;
           end 
          
      9'd481/*481:US*/:  begin 
           xpc10 <= 9'd482/*482:xpc10:482*/;
           A_SINT[19'h6_1fe8+11'h4d0] <= 32'd0;
           end 
          
      9'd482/*482:US*/:  begin 
           xpc10 <= 9'd483/*483:xpc10:483*/;
           A_SINT[19'h6_1fe8+11'h4d4] <= -32'd3;
           end 
          
      9'd483/*483:US*/:  begin 
           xpc10 <= 9'd484/*484:xpc10:484*/;
           A_SINT[19'h6_1fe8+11'h4d8] <= -32'd2;
           end 
          
      9'd484/*484:US*/:  begin 
           xpc10 <= 9'd485/*485:xpc10:485*/;
           A_SINT[19'h6_1fe8+11'h4dc] <= 32'd1;
           end 
          
      9'd485/*485:US*/:  begin 
           xpc10 <= 9'd486/*486:xpc10:486*/;
           A_SINT[19'h6_1fe8+11'h4e0] <= 32'd1;
           end 
          
      9'd486/*486:US*/:  begin 
           xpc10 <= 9'd487/*487:xpc10:487*/;
           A_SINT[19'h6_1fe8+11'h4e4] <= -32'd1;
           end 
          
      9'd487/*487:US*/:  begin 
           xpc10 <= 9'd488/*488:xpc10:488*/;
           A_SINT[19'h6_1fe8+11'h4e8] <= 32'd0;
           end 
          
      9'd488/*488:US*/:  begin 
           xpc10 <= 9'd489/*489:xpc10:489*/;
           A_SINT[19'h6_1fe8+11'h4ec] <= 32'd2;
           end 
          
      9'd489/*489:US*/:  begin 
           xpc10 <= 9'd490/*490:xpc10:490*/;
           A_SINT[19'h6_1fe8+11'h4f0] <= 32'd1;
           end 
          
      9'd490/*490:US*/:  begin 
           xpc10 <= 9'd491/*491:xpc10:491*/;
           A_SINT[19'h6_1fe8+11'h4f4] <= -32'd1;
           end 
          
      9'd491/*491:US*/:  begin 
           xpc10 <= 9'd492/*492:xpc10:492*/;
           A_SINT[19'h6_1fe8+11'h4f8] <= -32'd2;
           end 
          
      9'd492/*492:US*/:  begin 
           xpc10 <= 9'd493/*493:xpc10:493*/;
           A_SINT[19'h6_1fe8+11'h4fc] <= -32'd3;
           end 
          
      9'd493/*493:US*/:  begin 
           xpc10 <= 9'd494/*494:xpc10:494*/;
           A_SINT[19'h6_1fe8+11'h500] <= 32'd1;
           end 
          
      9'd494/*494:US*/:  begin 
           xpc10 <= 9'd495/*495:xpc10:495*/;
           A_SINT[19'h6_1fe8+11'h504] <= -32'd2;
           end 
          
      9'd495/*495:US*/:  begin 
           xpc10 <= 9'd496/*496:xpc10:496*/;
           A_SINT[19'h6_1fe8+11'h508] <= 32'd0;
           end 
          
      9'd496/*496:US*/:  begin 
           xpc10 <= 9'd497/*497:xpc10:497*/;
           A_SINT[19'h6_1fe8+11'h50c] <= 32'd0;
           end 
          
      9'd497/*497:US*/:  begin 
           xpc10 <= 9'd498/*498:xpc10:498*/;
           A_SINT[19'h6_1fe8+11'h510] <= -32'd3;
           end 
          
      9'd498/*498:US*/:  begin 
           xpc10 <= 9'd499/*499:xpc10:499*/;
           A_SINT[19'h6_1fe8+11'h514] <= 32'd0;
           end 
          
      9'd499/*499:US*/:  begin 
           xpc10 <= 9'd500/*500:xpc10:500*/;
           A_SINT[19'h6_1fe8+11'h518] <= -32'd1;
           end 
          
      9'd500/*500:US*/:  begin 
           xpc10 <= 9'd501/*501:xpc10:501*/;
           A_SINT[19'h6_1fe8+11'h51c] <= 32'd0;
           end 
          
      9'd501/*501:US*/:  begin 
           xpc10 <= 9'd502/*502:xpc10:502*/;
           A_SINT[19'h6_1fe8+11'h520] <= 32'd0;
           end 
          
      9'd502/*502:US*/:  begin 
           xpc10 <= 9'd503/*503:xpc10:503*/;
           A_SINT[19'h6_1fe8+11'h524] <= -32'd2;
           end 
          
      9'd503/*503:US*/:  begin 
           xpc10 <= 9'd504/*504:xpc10:504*/;
           A_SINT[19'h6_1fe8+11'h528] <= -32'd1;
           end 
          
      9'd504/*504:US*/:  begin 
           xpc10 <= 9'd505/*505:xpc10:505*/;
           A_SINT[19'h6_1fe8+11'h52c] <= 32'd0;
           end 
          
      9'd505/*505:US*/:  begin 
           xpc10 <= 9'd506/*506:xpc10:506*/;
           A_SINT[19'h6_1fe8+11'h530] <= 32'd0;
           end 
          
      9'd506/*506:US*/:  begin 
           xpc10 <= 9'd507/*507:xpc10:507*/;
           A_SINT[19'h6_1fe8+11'h534] <= -32'd1;
           end 
          
      9'd507/*507:US*/:  begin 
           xpc10 <= 9'd508/*508:xpc10:508*/;
           A_SINT[19'h6_1fe8+11'h538] <= -32'd1;
           end 
          
      9'd508/*508:US*/:  begin 
           xpc10 <= 9'd509/*509:xpc10:509*/;
           A_SINT[19'h6_1fe8+11'h53c] <= 32'd1;
           end 
          
      9'd509/*509:US*/:  begin 
           xpc10 <= 9'd510/*510:xpc10:510*/;
           A_SINT[19'h6_1fe8+11'h540] <= 32'd3;
           end 
          
      9'd510/*510:US*/:  begin 
           xpc10 <= 9'd511/*511:xpc10:511*/;
           A_SINT[19'h6_1fe8+11'h544] <= 32'd0;
           end 
          
      9'd511/*511:US*/:  begin 
           xpc10 <= 10'd512/*512:xpc10:512*/;
           A_SINT[19'h6_1fe8+11'h548] <= -32'd5;
           end 
          
      10'd512/*512:US*/:  begin 
           xpc10 <= 10'd513/*513:xpc10:513*/;
           A_SINT[19'h6_1fe8+11'h54c] <= -32'd3;
           end 
          
      10'd513/*513:US*/:  begin 
           xpc10 <= 10'd514/*514:xpc10:514*/;
           A_SINT[19'h6_1fe8+11'h550] <= 32'd0;
           end 
          
      10'd514/*514:US*/:  begin 
           xpc10 <= 10'd515/*515:xpc10:515*/;
           A_SINT[19'h6_1fe8+11'h554] <= -32'd2;
           end 
          
      10'd515/*515:US*/:  begin 
           xpc10 <= 10'd516/*516:xpc10:516*/;
           A_SINT[19'h6_1fe8+11'h558] <= -32'd2;
           end 
          
      10'd516/*516:US*/:  begin 
           xpc10 <= 10'd517/*517:xpc10:517*/;
           A_SINT[19'h6_1fe8+11'h55c] <= -32'd2;
           end 
          
      10'd517/*517:US*/:  begin 
           xpc10 <= 10'd518/*518:xpc10:518*/;
           A_SINT[19'h6_1fe8+11'h560] <= -32'd1;
           end 
          
      10'd518/*518:US*/:  begin 
           xpc10 <= 10'd519/*519:xpc10:519*/;
           A_SINT[19'h6_1fe8+11'h564] <= -32'd1;
           end 
          
      10'd519/*519:US*/:  begin 
           xpc10 <= 10'd520/*520:xpc10:520*/;
           A_SINT[19'h6_1fe8+11'h568] <= -32'd2;
           end 
          
      10'd520/*520:US*/:  begin 
           xpc10 <= 10'd521/*521:xpc10:521*/;
           A_SINT[19'h6_1fe8+11'h56c] <= 32'd4;
           end 
          
      10'd521/*521:US*/:  begin 
           xpc10 <= 10'd522/*522:xpc10:522*/;
           A_SINT[19'h6_1fe8+11'h570] <= -32'd2;
           end 
          
      10'd522/*522:US*/:  begin 
           xpc10 <= 10'd523/*523:xpc10:523*/;
           A_SINT[19'h6_1fe8+11'h574] <= 32'd2;
           end 
          
      10'd523/*523:US*/:  begin 
           xpc10 <= 10'd524/*524:xpc10:524*/;
           A_SINT[19'h6_1fe8+11'h578] <= 32'd2;
           end 
          
      10'd524/*524:US*/:  begin 
           xpc10 <= 10'd525/*525:xpc10:525*/;
           A_SINT[19'h6_1fe8+11'h57c] <= -32'd2;
           end 
          
      10'd525/*525:US*/:  begin 
           xpc10 <= 10'd526/*526:xpc10:526*/;
           A_SINT[19'h6_1fe8+11'h580] <= -32'd1;
           end 
          
      10'd526/*526:US*/:  begin 
           xpc10 <= 10'd527/*527:xpc10:527*/;
           A_SINT[19'h6_1fe8+11'h584] <= -32'd2;
           end 
          
      10'd527/*527:US*/:  begin 
           xpc10 <= 10'd528/*528:xpc10:528*/;
           A_SINT[19'h6_1fe8+11'h588] <= -32'd2;
           end 
          
      10'd528/*528:US*/:  begin 
           xpc10 <= 10'd529/*529:xpc10:529*/;
           A_SINT[19'h6_1fe8+11'h58c] <= -32'd1;
           end 
          
      10'd529/*529:US*/:  begin 
           xpc10 <= 10'd530/*530:xpc10:530*/;
           A_SINT[19'h6_1fe8+11'h590] <= 32'd0;
           end 
          
      10'd530/*530:US*/:  begin 
           xpc10 <= 10'd531/*531:xpc10:531*/;
           A_SINT[19'h6_1fe8+11'h594] <= 32'd4;
           end 
          
      10'd531/*531:US*/:  begin 
           xpc10 <= 10'd532/*532:xpc10:532*/;
           A_SINT[19'h6_1fe8+11'h598] <= -32'd6;
           end 
          
      10'd532/*532:US*/:  begin 
           xpc10 <= 10'd533/*533:xpc10:533*/;
           A_SINT[19'h6_1fe8+11'h59c] <= -32'd2;
           end 
          
      10'd533/*533:US*/:  begin 
           xpc10 <= 10'd534/*534:xpc10:534*/;
           A_SINT[19'h6_1fe8+11'h5a0] <= -32'd6;
           end 
          
      10'd534/*534:US*/:  begin 
           xpc10 <= 10'd535/*535:xpc10:535*/;
           A_SINT[19'h6_1fe8+11'h5a4] <= -32'd8;
           end 
          
      10'd535/*535:US*/:  begin 
           xpc10 <= 10'd536/*536:xpc10:536*/;
           A_SINT[19'h6_1fe8+11'h5a8] <= -32'd7;
           end 
          
      10'd536/*536:US*/:  begin 
           xpc10 <= 10'd537/*537:xpc10:537*/;
           A_SINT[19'h6_1fe8+11'h5ac] <= -32'd7;
           end 
          
      10'd537/*537:US*/:  begin 
           xpc10 <= 10'd538/*538:xpc10:538*/;
           A_SINT[19'h6_1fe8+11'h5b0] <= 32'd0;
           end 
          
      10'd538/*538:US*/:  begin 
           xpc10 <= 10'd539/*539:xpc10:539*/;
           A_SINT[19'h6_1fe8+11'h5b4] <= -32'd7;
           end 
          
      10'd539/*539:US*/:  begin 
           xpc10 <= 10'd540/*540:xpc10:540*/;
           A_SINT[19'h6_1fe8+11'h5b8] <= -32'd3;
           end 
          
      10'd540/*540:US*/:  begin 
           xpc10 <= 10'd541/*541:xpc10:541*/;
           A_SINT[19'h6_1fe8+11'h5bc] <= -32'd5;
           end 
          
      10'd541/*541:US*/:  begin 
           xpc10 <= 10'd542/*542:xpc10:542*/;
           A_SINT[19'h6_1fe8+11'h5c0] <= -32'd3;
           end 
          
      10'd542/*542:US*/:  begin 
           xpc10 <= 10'd543/*543:xpc10:543*/;
           A_SINT[19'h6_1fe8+11'h5c4] <= -32'd2;
           end 
          
      10'd543/*543:US*/:  begin 
           xpc10 <= 10'd544/*544:xpc10:544*/;
           A_SINT[19'h6_1fe8+11'h5c8] <= -32'd4;
           end 
          
      10'd544/*544:US*/:  begin 
           xpc10 <= 10'd545/*545:xpc10:545*/;
           A_SINT[19'h6_1fe8+11'h5cc] <= -32'd4;
           end 
          
      10'd545/*545:US*/:  begin 
           xpc10 <= 10'd546/*546:xpc10:546*/;
           A_SINT[19'h6_1fe8+11'h5d0] <= -32'd6;
           end 
          
      10'd546/*546:US*/:  begin 
           xpc10 <= 10'd547/*547:xpc10:547*/;
           A_SINT[19'h6_1fe8+11'h5d4] <= -32'd5;
           end 
          
      10'd547/*547:US*/:  begin 
           xpc10 <= 10'd548/*548:xpc10:548*/;
           A_SINT[19'h6_1fe8+11'h5d8] <= 32'd2;
           end 
          
      10'd548/*548:US*/:  begin 
           xpc10 <= 10'd549/*549:xpc10:549*/;
           A_SINT[19'h6_1fe8+11'h5dc] <= -32'd2;
           end 
          
      10'd549/*549:US*/:  begin 
           xpc10 <= 10'd550/*550:xpc10:550*/;
           A_SINT[19'h6_1fe8+11'h5e0] <= -32'd5;
           end 
          
      10'd550/*550:US*/:  begin 
           xpc10 <= 10'd551/*551:xpc10:551*/;
           A_SINT[19'h6_1fe8+11'h5e4] <= -32'd6;
           end 
          
      10'd551/*551:US*/:  begin 
           xpc10 <= 10'd552/*552:xpc10:552*/;
           A_SINT[19'h6_1fe8+11'h5e8] <= 32'd17;
           end 
          
      10'd552/*552:US*/:  begin 
           xpc10 <= 10'd553/*553:xpc10:553*/;
           A_SINT[19'h6_1fe8+11'h5ec] <= 32'd0;
           end 
          
      10'd553/*553:US*/:  begin 
           xpc10 <= 10'd554/*554:xpc10:554*/;
           A_SINT[19'h6_1fe8+11'h5f0] <= -32'd3;
           end 
          
      10'd554/*554:US*/:  begin 
           xpc10 <= 10'd555/*555:xpc10:555*/;
           A_SINT[19'h6_1fe8+11'h5f4] <= 32'd0;
           end 
          
      10'd555/*555:US*/:  begin 
           xpc10 <= 10'd556/*556:xpc10:556*/;
           A_SINT[19'h6_1fe8+11'h5f8] <= -32'd4;
           end 
          
      10'd556/*556:US*/:  begin 
           xpc10 <= 10'd557/*557:xpc10:557*/;
           A_SINT[19'h6_1fe8+11'h5fc] <= -32'd4;
           end 
          
      10'd557/*557:US*/:  begin 
           xpc10 <= 10'd558/*558:xpc10:558*/;
           A_SINT[19'h6_1fe8+11'h600] <= 32'd7;
           end 
          
      10'd558/*558:US*/:  begin 
           xpc10 <= 10'd559/*559:xpc10:559*/;
           A_SINT[19'h6_1fe8+11'h604] <= -32'd5;
           end 
          
      10'd559/*559:US*/:  begin 
           xpc10 <= 10'd560/*560:xpc10:560*/;
           A_SINT[19'h6_1fe8+11'h608] <= 32'd0;
           end 
          
      10'd560/*560:US*/:  begin 
           xpc10 <= 10'd561/*561:xpc10:561*/;
           A_SINT[19'h6_1fe8+11'h60c] <= -32'd1;
           end 
          
      10'd561/*561:US*/:  begin 
           xpc10 <= 10'd562/*562:xpc10:562*/;
           A_SINT[19'h6_1fe8+11'h610] <= -32'd4;
           end 
          
      10'd562/*562:US*/:  begin 
           xpc10 <= 10'd563/*563:xpc10:563*/;
           A_SINT[19'h6_1fe8+11'h614] <= -32'd1;
           end 
          
      10'd563/*563:US*/:  begin 
           xpc10 <= 10'd564/*564:xpc10:564*/;
           A_SINT[19'h6_1fe8+11'h618] <= -32'd2;
           end 
          
      10'd564/*564:US*/:  begin 
           xpc10 <= 10'd565/*565:xpc10:565*/;
           A_SINT[19'h6_1fe8+11'h61c] <= -32'd2;
           end 
          
      10'd565/*565:US*/:  begin 
           xpc10 <= 10'd566/*566:xpc10:566*/;
           A_SINT[19'h6_1fe8+11'h620] <= -32'd5;
           end 
          
      10'd566/*566:US*/:  begin 
           xpc10 <= 10'd567/*567:xpc10:567*/;
           A_SINT[19'h6_1fe8+11'h624] <= -32'd4;
           end 
          
      10'd567/*567:US*/:  begin 
           xpc10 <= 10'd568/*568:xpc10:568*/;
           A_SINT[19'h6_1fe8+11'h628] <= -32'd4;
           end 
          
      10'd568/*568:US*/:  begin 
           xpc10 <= 10'd569/*569:xpc10:569*/;
           A_SINT[19'h6_1fe8+11'h62c] <= -32'd3;
           end 
          
      10'd569/*569:US*/:  begin 
           xpc10 <= 10'd570/*570:xpc10:570*/;
           A_SINT[19'h6_1fe8+11'h630] <= -32'd3;
           end 
          
      10'd570/*570:US*/:  begin 
           xpc10 <= 10'd571/*571:xpc10:571*/;
           A_SINT[19'h6_1fe8+11'h634] <= -32'd2;
           end 
          
      10'd571/*571:US*/:  begin 
           xpc10 <= 10'd572/*572:xpc10:572*/;
           A_SINT[19'h6_1fe8+11'h638] <= 32'd0;
           end 
          
      10'd572/*572:US*/:  begin 
           xpc10 <= 10'd573/*573:xpc10:573*/;
           A_UINT[19'h6_1a80+0] <= 32'd0;
           A_SINT[19'h6_1fe8+11'h63c] <= 32'd10;
           end 
          
      10'd573/*573:US*/:  begin 
           xpc10 <= 10'd574/*574:xpc10:574*/;
           A_UINT[19'h6_1a80+3'h4] <= 32'd79764919;
           end 
          
      10'd574/*574:US*/:  begin 
           xpc10 <= 10'd575/*575:xpc10:575*/;
           A_UINT[19'h6_1a80+4'h8] <= 32'd159529838;
           end 
          
      10'd575/*575:US*/:  begin 
           xpc10 <= 10'd576/*576:xpc10:576*/;
           A_UINT[19'h6_1a80+4'hc] <= 32'd222504665;
           end 
          
      10'd576/*576:US*/:  begin 
           xpc10 <= 10'd577/*577:xpc10:577*/;
           A_UINT[19'h6_1a80+5'h10] <= 32'd319059676;
           end 
          
      10'd577/*577:US*/:  begin 
           xpc10 <= 10'd578/*578:xpc10:578*/;
           A_UINT[19'h6_1a80+5'h14] <= 32'd398814059;
           end 
          
      10'd578/*578:US*/:  begin 
           xpc10 <= 10'd579/*579:xpc10:579*/;
           A_UINT[19'h6_1a80+5'h18] <= 32'd445009330;
           end 
          
      10'd579/*579:US*/:  begin 
           xpc10 <= 10'd580/*580:xpc10:580*/;
           A_UINT[19'h6_1a80+5'h1c] <= 32'd507990021;
           end 
          
      10'd580/*580:US*/:  begin 
           xpc10 <= 10'd581/*581:xpc10:581*/;
           A_UINT[19'h6_1a80+6'h20] <= 32'd638119352;
           end 
          
      10'd581/*581:US*/:  begin 
           xpc10 <= 10'd582/*582:xpc10:582*/;
           A_UINT[19'h6_1a80+6'h24] <= 32'd583659535;
           end 
          
      10'd582/*582:US*/:  begin 
           xpc10 <= 10'd583/*583:xpc10:583*/;
           A_UINT[19'h6_1a80+6'h28] <= 32'd797628118;
           end 
          
      10'd583/*583:US*/:  begin 
           xpc10 <= 10'd584/*584:xpc10:584*/;
           A_UINT[19'h6_1a80+6'h2c] <= 32'd726387553;
           end 
          
      10'd584/*584:US*/:  begin 
           xpc10 <= 10'd585/*585:xpc10:585*/;
           A_UINT[19'h6_1a80+6'h30] <= 32'd890018660;
           end 
          
      10'd585/*585:US*/:  begin 
           xpc10 <= 10'd586/*586:xpc10:586*/;
           A_UINT[19'h6_1a80+6'h34] <= 32'd835552979;
           end 
          
      10'd586/*586:US*/:  begin 
           xpc10 <= 10'd587/*587:xpc10:587*/;
           A_UINT[19'h6_1a80+6'h38] <= 32'd1015980042;
           end 
          
      10'd587/*587:US*/:  begin 
           xpc10 <= 10'd588/*588:xpc10:588*/;
           A_UINT[19'h6_1a80+6'h3c] <= 32'd944750013;
           end 
          
      10'd588/*588:US*/:  begin 
           xpc10 <= 10'd589/*589:xpc10:589*/;
           A_UINT[19'h6_1a80+7'h40] <= 32'd1276238704;
           end 
          
      10'd589/*589:US*/:  begin 
           xpc10 <= 10'd590/*590:xpc10:590*/;
           A_UINT[19'h6_1a80+7'h44] <= 32'd1221641927;
           end 
          
      10'd590/*590:US*/:  begin 
           xpc10 <= 10'd591/*591:xpc10:591*/;
           A_UINT[19'h6_1a80+7'h48] <= 32'd1167319070;
           end 
          
      10'd591/*591:US*/:  begin 
           xpc10 <= 10'd592/*592:xpc10:592*/;
           A_UINT[19'h6_1a80+7'h4c] <= 32'd1095957929;
           end 
          
      10'd592/*592:US*/:  begin 
           xpc10 <= 10'd593/*593:xpc10:593*/;
           A_UINT[19'h6_1a80+7'h50] <= 32'd1595256236;
           end 
          
      10'd593/*593:US*/:  begin 
           xpc10 <= 10'd594/*594:xpc10:594*/;
           A_UINT[19'h6_1a80+7'h54] <= 32'd1540665371;
           end 
          
      10'd594/*594:US*/:  begin 
           xpc10 <= 10'd595/*595:xpc10:595*/;
           A_UINT[19'h6_1a80+7'h58] <= 32'd1452775106;
           end 
          
      10'd595/*595:US*/:  begin 
           xpc10 <= 10'd596/*596:xpc10:596*/;
           A_UINT[19'h6_1a80+7'h5c] <= 32'd1381403509;
           end 
          
      10'd596/*596:US*/:  begin 
           xpc10 <= 10'd597/*597:xpc10:597*/;
           A_UINT[19'h6_1a80+7'h60] <= 32'd1780037320;
           end 
          
      10'd597/*597:US*/:  begin 
           xpc10 <= 10'd598/*598:xpc10:598*/;
           A_UINT[19'h6_1a80+7'h64] <= 32'd1859660671;
           end 
          
      10'd598/*598:US*/:  begin 
           xpc10 <= 10'd599/*599:xpc10:599*/;
           A_UINT[19'h6_1a80+7'h68] <= 32'd1671105958;
           end 
          
      10'd599/*599:US*/:  begin 
           xpc10 <= 10'd600/*600:xpc10:600*/;
           A_UINT[19'h6_1a80+7'h6c] <= 32'd1733955601;
           end 
          
      10'd600/*600:US*/:  begin 
           xpc10 <= 10'd601/*601:xpc10:601*/;
           A_UINT[19'h6_1a80+7'h70] <= 32'd2031960084;
           end 
          
      10'd601/*601:US*/:  begin 
           xpc10 <= 10'd602/*602:xpc10:602*/;
           A_UINT[19'h6_1a80+7'h74] <= 32'd2111593891;
           end 
          
      10'd602/*602:US*/:  begin 
           xpc10 <= 10'd603/*603:xpc10:603*/;
           A_UINT[19'h6_1a80+7'h78] <= 32'd1889500026;
           end 
          
      10'd603/*603:US*/:  begin 
           xpc10 <= 10'd604/*604:xpc10:604*/;
           A_UINT[19'h6_1a80+7'h7c] <= 32'd1952343757;
           end 
          
      10'd604/*604:US*/:  begin 
           xpc10 <= 10'd605/*605:xpc10:605*/;
           A_UINT[19'h6_1a80+8'h80] <= -32'd1742489888;
           end 
          
      10'd605/*605:US*/:  begin 
           xpc10 <= 10'd606/*606:xpc10:606*/;
           A_UINT[19'h6_1a80+8'h84] <= -32'd1662866601;
           end 
          
      10'd606/*606:US*/:  begin 
           xpc10 <= 10'd607/*607:xpc10:607*/;
           A_UINT[19'h6_1a80+8'h88] <= -32'd1851683442;
           end 
          
      10'd607/*607:US*/:  begin 
           xpc10 <= 10'd608/*608:xpc10:608*/;
           A_UINT[19'h6_1a80+8'h8c] <= -32'd1788833735;
           end 
          
      10'd608/*608:US*/:  begin 
           xpc10 <= 10'd609/*609:xpc10:609*/;
           A_UINT[19'h6_1a80+8'h90] <= -32'd1960329156;
           end 
          
      10'd609/*609:US*/:  begin 
           xpc10 <= 10'd610/*610:xpc10:610*/;
           A_UINT[19'h6_1a80+8'h94] <= -32'd1880695413;
           end 
          
      10'd610/*610:US*/:  begin 
           xpc10 <= 10'd611/*611:xpc10:611*/;
           A_UINT[19'h6_1a80+8'h98] <= -32'd2103051438;
           end 
          
      10'd611/*611:US*/:  begin 
           xpc10 <= 10'd612/*612:xpc10:612*/;
           A_UINT[19'h6_1a80+8'h9c] <= -32'd2040207643;
           end 
          
      10'd612/*612:US*/:  begin 
           xpc10 <= 10'd613/*613:xpc10:613*/;
           A_UINT[19'h6_1a80+8'ha0] <= -32'd1104454824;
           end 
          
      10'd613/*613:US*/:  begin 
           xpc10 <= 10'd614/*614:xpc10:614*/;
           A_UINT[19'h6_1a80+8'ha4] <= -32'd1159051537;
           end 
          
      10'd614/*614:US*/:  begin 
           xpc10 <= 10'd615/*615:xpc10:615*/;
           A_UINT[19'h6_1a80+8'ha8] <= -32'd1213636554;
           end 
          
      10'd615/*615:US*/:  begin 
           xpc10 <= 10'd616/*616:xpc10:616*/;
           A_UINT[19'h6_1a80+8'hac] <= -32'd1284997759;
           end 
          
      10'd616/*616:US*/:  begin 
           xpc10 <= 10'd617/*617:xpc10:617*/;
           A_UINT[19'h6_1a80+8'hb0] <= -32'd1389417084;
           end 
          
      10'd617/*617:US*/:  begin 
           xpc10 <= 10'd618/*618:xpc10:618*/;
           A_UINT[19'h6_1a80+8'hb4] <= -32'd1444007885;
           end 
          
      10'd618/*618:US*/:  begin 
           xpc10 <= 10'd619/*619:xpc10:619*/;
           A_UINT[19'h6_1a80+8'hb8] <= -32'd1532160278;
           end 
          
      10'd619/*619:US*/:  begin 
           xpc10 <= 10'd620/*620:xpc10:620*/;
           A_UINT[19'h6_1a80+8'hbc] <= -32'd1603531939;
           end 
          
      10'd620/*620:US*/:  begin 
           xpc10 <= 10'd621/*621:xpc10:621*/;
           A_UINT[19'h6_1a80+8'hc0] <= -32'd734892656;
           end 
          
      10'd621/*621:US*/:  begin 
           xpc10 <= 10'd622/*622:xpc10:622*/;
           A_UINT[19'h6_1a80+8'hc4] <= -32'd789352409;
           end 
          
      10'd622/*622:US*/:  begin 
           xpc10 <= 10'd623/*623:xpc10:623*/;
           A_UINT[19'h6_1a80+8'hc8] <= -32'd575645954;
           end 
          
      10'd623/*623:US*/:  begin 
           xpc10 <= 10'd624/*624:xpc10:624*/;
           A_UINT[19'h6_1a80+8'hcc] <= -32'd646886583;
           end 
          
      10'd624/*624:US*/:  begin 
           xpc10 <= 10'd625/*625:xpc10:625*/;
           A_UINT[19'h6_1a80+8'hd0] <= -32'd952755380;
           end 
          
      10'd625/*625:US*/:  begin 
           xpc10 <= 10'd626/*626:xpc10:626*/;
           A_UINT[19'h6_1a80+8'hd4] <= -32'd1007220997;
           end 
          
      10'd626/*626:US*/:  begin 
           xpc10 <= 10'd627/*627:xpc10:627*/;
           A_UINT[19'h6_1a80+8'hd8] <= -32'd827056094;
           end 
          
      10'd627/*627:US*/:  begin 
           xpc10 <= 10'd628/*628:xpc10:628*/;
           A_UINT[19'h6_1a80+8'hdc] <= -32'd898286187;
           end 
          
      10'd628/*628:US*/:  begin 
           xpc10 <= 10'd629/*629:xpc10:629*/;
           A_UINT[19'h6_1a80+8'he0] <= -32'd231047128;
           end 
          
      10'd629/*629:US*/:  begin 
           xpc10 <= 10'd630/*630:xpc10:630*/;
           A_UINT[19'h6_1a80+8'he4] <= -32'd151282273;
           end 
          
      10'd630/*630:US*/:  begin 
           xpc10 <= 10'd631/*631:xpc10:631*/;
           A_UINT[19'h6_1a80+8'he8] <= -32'd71779514;
           end 
          
      10'd631/*631:US*/:  begin 
           xpc10 <= 10'd632/*632:xpc10:632*/;
           A_UINT[19'h6_1a80+8'hec] <= -32'd8804623;
           end 
          
      10'd632/*632:US*/:  begin 
           xpc10 <= 10'd633/*633:xpc10:633*/;
           A_UINT[19'h6_1a80+8'hf0] <= -32'd515967244;
           end 
          
      10'd633/*633:US*/:  begin 
           xpc10 <= 10'd634/*634:xpc10:634*/;
           A_UINT[19'h6_1a80+8'hf4] <= -32'd436212925;
           end 
          
      10'd634/*634:US*/:  begin 
           xpc10 <= 10'd635/*635:xpc10:635*/;
           A_UINT[19'h6_1a80+8'hf8] <= -32'd390279782;
           end 
          
      10'd635/*635:US*/:  begin 
           xpc10 <= 10'd636/*636:xpc10:636*/;
           A_UINT[19'h6_1a80+8'hfc] <= -32'd327299027;
           end 
          
      10'd636/*636:US*/:  begin 
           xpc10 <= 10'd637/*637:xpc10:637*/;
           A_UINT[19'h6_1a80+9'h100] <= 32'd881225847;
           end 
          
      10'd637/*637:US*/:  begin 
           xpc10 <= 10'd638/*638:xpc10:638*/;
           A_UINT[19'h6_1a80+9'h104] <= 32'd809987520;
           end 
          
      10'd638/*638:US*/:  begin 
           xpc10 <= 10'd639/*639:xpc10:639*/;
           A_UINT[19'h6_1a80+9'h108] <= 32'd1023691545;
           end 
          
      10'd639/*639:US*/:  begin 
           xpc10 <= 10'd640/*640:xpc10:640*/;
           A_UINT[19'h6_1a80+9'h10c] <= 32'd969234094;
           end 
          
      10'd640/*640:US*/:  begin 
           xpc10 <= 10'd641/*641:xpc10:641*/;
           A_UINT[19'h6_1a80+9'h110] <= 32'd662832811;
           end 
          
      10'd641/*641:US*/:  begin 
           xpc10 <= 10'd642/*642:xpc10:642*/;
           A_UINT[19'h6_1a80+9'h114] <= 32'd591600412;
           end 
          
      10'd642/*642:US*/:  begin 
           xpc10 <= 10'd643/*643:xpc10:643*/;
           A_UINT[19'h6_1a80+9'h118] <= 32'd771767749;
           end 
          
      10'd643/*643:US*/:  begin 
           xpc10 <= 10'd644/*644:xpc10:644*/;
           A_UINT[19'h6_1a80+9'h11c] <= 32'd717299826;
           end 
          
      10'd644/*644:US*/:  begin 
           xpc10 <= 10'd645/*645:xpc10:645*/;
           A_UINT[19'h6_1a80+9'h120] <= 32'd311336399;
           end 
          
      10'd645/*645:US*/:  begin 
           xpc10 <= 10'd646/*646:xpc10:646*/;
           A_UINT[19'h6_1a80+9'h124] <= 32'd374308984;
           end 
          
      10'd646/*646:US*/:  begin 
           xpc10 <= 10'd647/*647:xpc10:647*/;
           A_UINT[19'h6_1a80+9'h128] <= 32'd453813921;
           end 
          
      10'd647/*647:US*/:  begin 
           xpc10 <= 10'd648/*648:xpc10:648*/;
           A_UINT[19'h6_1a80+9'h12c] <= 32'd533576470;
           end 
          
      10'd648/*648:US*/:  begin 
           xpc10 <= 10'd649/*649:xpc10:649*/;
           A_UINT[19'h6_1a80+9'h130] <= 32'd25881363;
           end 
          
      10'd649/*649:US*/:  begin 
           xpc10 <= 10'd650/*650:xpc10:650*/;
           A_UINT[19'h6_1a80+9'h134] <= 32'd88864420;
           end 
          
      10'd650/*650:US*/:  begin 
           xpc10 <= 10'd651/*651:xpc10:651*/;
           A_UINT[19'h6_1a80+9'h138] <= 32'd134795389;
           end 
          
      10'd651/*651:US*/:  begin 
           xpc10 <= 10'd652/*652:xpc10:652*/;
           A_UINT[19'h6_1a80+9'h13c] <= 32'd214552010;
           end 
          
      10'd652/*652:US*/:  begin 
           xpc10 <= 10'd653/*653:xpc10:653*/;
           A_UINT[19'h6_1a80+9'h140] <= 32'd2023205639;
           end 
          
      10'd653/*653:US*/:  begin 
           xpc10 <= 10'd654/*654:xpc10:654*/;
           A_UINT[19'h6_1a80+9'h144] <= 32'd2086057648;
           end 
          
      10'd654/*654:US*/:  begin 
           xpc10 <= 10'd655/*655:xpc10:655*/;
           A_UINT[19'h6_1a80+9'h148] <= 32'd1897238633;
           end 
          
      10'd655/*655:US*/:  begin 
           xpc10 <= 10'd656/*656:xpc10:656*/;
           A_UINT[19'h6_1a80+9'h14c] <= 32'd1976864222;
           end 
          
      10'd656/*656:US*/:  begin 
           xpc10 <= 10'd657/*657:xpc10:657*/;
           A_UINT[19'h6_1a80+9'h150] <= 32'd1804852699;
           end 
          
      10'd657/*657:US*/:  begin 
           xpc10 <= 10'd658/*658:xpc10:658*/;
           A_UINT[19'h6_1a80+9'h154] <= 32'd1867694188;
           end 
          
      10'd658/*658:US*/:  begin 
           xpc10 <= 10'd659/*659:xpc10:659*/;
           A_UINT[19'h6_1a80+9'h158] <= 32'd1645340341;
           end 
          
      10'd659/*659:US*/:  begin 
           xpc10 <= 10'd660/*660:xpc10:660*/;
           A_UINT[19'h6_1a80+9'h15c] <= 32'd1724971778;
           end 
          
      10'd660/*660:US*/:  begin 
           xpc10 <= 10'd661/*661:xpc10:661*/;
           A_UINT[19'h6_1a80+9'h160] <= 32'd1587496639;
           end 
          
      10'd661/*661:US*/:  begin 
           xpc10 <= 10'd662/*662:xpc10:662*/;
           A_UINT[19'h6_1a80+9'h164] <= 32'd1516133128;
           end 
          
      10'd662/*662:US*/:  begin 
           xpc10 <= 10'd663/*663:xpc10:663*/;
           A_UINT[19'h6_1a80+9'h168] <= 32'd1461550545;
           end 
          
      10'd663/*663:US*/:  begin 
           xpc10 <= 10'd664/*664:xpc10:664*/;
           A_UINT[19'h6_1a80+9'h16c] <= 32'd1406951526;
           end 
          
      10'd664/*664:US*/:  begin 
           xpc10 <= 10'd665/*665:xpc10:665*/;
           A_UINT[19'h6_1a80+9'h170] <= 32'd1302016099;
           end 
          
      10'd665/*665:US*/:  begin 
           xpc10 <= 10'd666/*666:xpc10:666*/;
           A_UINT[19'h6_1a80+9'h174] <= 32'd1230646740;
           end 
          
      10'd666/*666:US*/:  begin 
           xpc10 <= 10'd667/*667:xpc10:667*/;
           A_UINT[19'h6_1a80+9'h178] <= 32'd1142491917;
           end 
          
      10'd667/*667:US*/:  begin 
           xpc10 <= 10'd668/*668:xpc10:668*/;
           A_UINT[19'h6_1a80+9'h17c] <= 32'd1087903418;
           end 
          
      10'd668/*668:US*/:  begin 
           xpc10 <= 10'd669/*669:xpc10:669*/;
           A_UINT[19'h6_1a80+9'h180] <= -32'd1398421865;
           end 
          
      10'd669/*669:US*/:  begin 
           xpc10 <= 10'd670/*670:xpc10:670*/;
           A_UINT[19'h6_1a80+9'h184] <= -32'd1469785312;
           end 
          
      10'd670/*670:US*/:  begin 
           xpc10 <= 10'd671/*671:xpc10:671*/;
           A_UINT[19'h6_1a80+9'h188] <= -32'd1524105735;
           end 
          
      10'd671/*671:US*/:  begin 
           xpc10 <= 10'd672/*672:xpc10:672*/;
           A_UINT[19'h6_1a80+9'h18c] <= -32'd1578704818;
           end 
          
      10'd672/*672:US*/:  begin 
           xpc10 <= 10'd673/*673:xpc10:673*/;
           A_UINT[19'h6_1a80+9'h190] <= -32'd1079922613;
           end 
          
      10'd673/*673:US*/:  begin 
           xpc10 <= 10'd674/*674:xpc10:674*/;
           A_UINT[19'h6_1a80+9'h194] <= -32'd1151291908;
           end 
          
      10'd674/*674:US*/:  begin 
           xpc10 <= 10'd675/*675:xpc10:675*/;
           A_UINT[19'h6_1a80+9'h198] <= -32'd1239184603;
           end 
          
      10'd675/*675:US*/:  begin 
           xpc10 <= 10'd676/*676:xpc10:676*/;
           A_UINT[19'h6_1a80+9'h19c] <= -32'd1293773166;
           end 
          
      10'd676/*676:US*/:  begin 
           xpc10 <= 10'd677/*677:xpc10:677*/;
           A_UINT[19'h6_1a80+9'h1a0] <= -32'd1968362705;
           end 
          
      10'd677/*677:US*/:  begin 
           xpc10 <= 10'd678/*678:xpc10:678*/;
           A_UINT[19'h6_1a80+9'h1a4] <= -32'd1905510760;
           end 
          
      10'd678/*678:US*/:  begin 
           xpc10 <= 10'd679/*679:xpc10:679*/;
           A_UINT[19'h6_1a80+9'h1a8] <= -32'd2094067647;
           end 
          
      10'd679/*679:US*/:  begin 
           xpc10 <= 10'd680/*680:xpc10:680*/;
           A_UINT[19'h6_1a80+9'h1ac] <= -32'd2014441994;
           end 
          
      10'd680/*680:US*/:  begin 
           xpc10 <= 10'd681/*681:xpc10:681*/;
           A_UINT[19'h6_1a80+9'h1b0] <= -32'd1716953613;
           end 
          
      10'd681/*681:US*/:  begin 
           xpc10 <= 10'd682/*682:xpc10:682*/;
           A_UINT[19'h6_1a80+9'h1b4] <= -32'd1654112188;
           end 
          
      10'd682/*682:US*/:  begin 
           xpc10 <= 10'd683/*683:xpc10:683*/;
           A_UINT[19'h6_1a80+9'h1b8] <= -32'd1876203875;
           end 
          
      10'd683/*683:US*/:  begin 
           xpc10 <= 10'd684/*684:xpc10:684*/;
           A_UINT[19'h6_1a80+9'h1bc] <= -32'd1796572374;
           end 
          
      10'd684/*684:US*/:  begin 
           xpc10 <= 10'd685/*685:xpc10:685*/;
           A_UINT[19'h6_1a80+9'h1c0] <= -32'd525066777;
           end 
          
      10'd685/*685:US*/:  begin 
           xpc10 <= 10'd686/*686:xpc10:686*/;
           A_UINT[19'h6_1a80+9'h1c4] <= -32'd462094256;
           end 
          
      10'd686/*686:US*/:  begin 
           xpc10 <= 10'd687/*687:xpc10:687*/;
           A_UINT[19'h6_1a80+9'h1c8] <= -32'd382327159;
           end 
          
      10'd687/*687:US*/:  begin 
           xpc10 <= 10'd688/*688:xpc10:688*/;
           A_UINT[19'h6_1a80+9'h1cc] <= -32'd302564546;
           end 
          
      10'd688/*688:US*/:  begin 
           xpc10 <= 10'd689/*689:xpc10:689*/;
           A_UINT[19'h6_1a80+9'h1d0] <= -32'd206542021;
           end 
          
      10'd689/*689:US*/:  begin 
           xpc10 <= 10'd690/*690:xpc10:690*/;
           A_UINT[19'h6_1a80+9'h1d4] <= -32'd143559028;
           end 
          
      10'd690/*690:US*/:  begin 
           xpc10 <= 10'd691/*691:xpc10:691*/;
           A_UINT[19'h6_1a80+9'h1d8] <= -32'd97365931;
           end 
          
      10'd691/*691:US*/:  begin 
           xpc10 <= 10'd692/*692:xpc10:692*/;
           A_UINT[19'h6_1a80+9'h1dc] <= -32'd17609246;
           end 
          
      10'd692/*692:US*/:  begin 
           xpc10 <= 10'd693/*693:xpc10:693*/;
           A_UINT[19'h6_1a80+9'h1e0] <= -32'd960696225;
           end 
          
      10'd693/*693:US*/:  begin 
           xpc10 <= 10'd694/*694:xpc10:694*/;
           A_UINT[19'h6_1a80+9'h1e4] <= -32'd1031934488;
           end 
          
      10'd694/*694:US*/:  begin 
           xpc10 <= 10'd695/*695:xpc10:695*/;
           A_UINT[19'h6_1a80+9'h1e8] <= -32'd817968335;
           end 
          
      10'd695/*695:US*/:  begin 
           xpc10 <= 10'd696/*696:xpc10:696*/;
           A_UINT[19'h6_1a80+9'h1ec] <= -32'd872425850;
           end 
          
      10'd696/*696:US*/:  begin 
           xpc10 <= 10'd697/*697:xpc10:697*/;
           A_UINT[19'h6_1a80+9'h1f0] <= -32'd709327229;
           end 
          
      10'd697/*697:US*/:  begin 
           xpc10 <= 10'd698/*698:xpc10:698*/;
           A_UINT[19'h6_1a80+9'h1f4] <= -32'd780559564;
           end 
          
      10'd698/*698:US*/:  begin 
           xpc10 <= 10'd699/*699:xpc10:699*/;
           A_UINT[19'h6_1a80+9'h1f8] <= -32'd600130067;
           end 
          
      10'd699/*699:US*/:  begin 
           xpc10 <= 10'd700/*700:xpc10:700*/;
           A_UINT[19'h6_1a80+9'h1fc] <= -32'd654598054;
           end 
          
      10'd700/*700:US*/:  begin 
           xpc10 <= 10'd701/*701:xpc10:701*/;
           A_UINT[19'h6_1a80+10'h200] <= 32'd1762451694;
           end 
          
      10'd701/*701:US*/:  begin 
           xpc10 <= 10'd702/*702:xpc10:702*/;
           A_UINT[19'h6_1a80+10'h204] <= 32'd1842216281;
           end 
          
      10'd702/*702:US*/:  begin 
           xpc10 <= 10'd703/*703:xpc10:703*/;
           A_UINT[19'h6_1a80+10'h208] <= 32'd1619975040;
           end 
          
      10'd703/*703:US*/:  begin 
           xpc10 <= 10'd704/*704:xpc10:704*/;
           A_UINT[19'h6_1a80+10'h20c] <= 32'd1682949687;
           end 
          
      10'd704/*704:US*/:  begin 
           xpc10 <= 10'd705/*705:xpc10:705*/;
           A_UINT[19'h6_1a80+10'h210] <= 32'd2047383090;
           end 
          
      10'd705/*705:US*/:  begin 
           xpc10 <= 10'd706/*706:xpc10:706*/;
           A_UINT[19'h6_1a80+10'h214] <= 32'd2127137669;
           end 
          
      10'd706/*706:US*/:  begin 
           xpc10 <= 10'd707/*707:xpc10:707*/;
           A_UINT[19'h6_1a80+10'h218] <= 32'd1938468188;
           end 
          
      10'd707/*707:US*/:  begin 
           xpc10 <= 10'd708/*708:xpc10:708*/;
           A_UINT[19'h6_1a80+10'h21c] <= 32'd2001449195;
           end 
          
      10'd708/*708:US*/:  begin 
           xpc10 <= 10'd709/*709:xpc10:709*/;
           A_UINT[19'h6_1a80+10'h220] <= 32'd1325665622;
           end 
          
      10'd709/*709:US*/:  begin 
           xpc10 <= 10'd710/*710:xpc10:710*/;
           A_UINT[19'h6_1a80+10'h224] <= 32'd1271206113;
           end 
          
      10'd710/*710:US*/:  begin 
           xpc10 <= 10'd711/*711:xpc10:711*/;
           A_UINT[19'h6_1a80+10'h228] <= 32'd1183200824;
           end 
          
      10'd711/*711:US*/:  begin 
           xpc10 <= 10'd712/*712:xpc10:712*/;
           A_UINT[19'h6_1a80+10'h22c] <= 32'd1111960463;
           end 
          
      10'd712/*712:US*/:  begin 
           xpc10 <= 10'd713/*713:xpc10:713*/;
           A_UINT[19'h6_1a80+10'h230] <= 32'd1543535498;
           end 
          
      10'd713/*713:US*/:  begin 
           xpc10 <= 10'd714/*714:xpc10:714*/;
           A_UINT[19'h6_1a80+10'h234] <= 32'd1489069629;
           end 
          
      10'd714/*714:US*/:  begin 
           xpc10 <= 10'd715/*715:xpc10:715*/;
           A_UINT[19'h6_1a80+10'h238] <= 32'd1434599652;
           end 
          
      10'd715/*715:US*/:  begin 
           xpc10 <= 10'd716/*716:xpc10:716*/;
           A_UINT[19'h6_1a80+10'h23c] <= 32'd1363369299;
           end 
          
      10'd716/*716:US*/:  begin 
           xpc10 <= 10'd717/*717:xpc10:717*/;
           A_UINT[19'h6_1a80+10'h240] <= 32'd622672798;
           end 
          
      10'd717/*717:US*/:  begin 
           xpc10 <= 10'd718/*718:xpc10:718*/;
           A_UINT[19'h6_1a80+10'h244] <= 32'd568075817;
           end 
          
      10'd718/*718:US*/:  begin 
           xpc10 <= 10'd719/*719:xpc10:719*/;
           A_UINT[19'h6_1a80+10'h248] <= 32'd748617968;
           end 
          
      10'd719/*719:US*/:  begin 
           xpc10 <= 10'd720/*720:xpc10:720*/;
           A_UINT[19'h6_1a80+10'h24c] <= 32'd677256519;
           end 
          
      10'd720/*720:US*/:  begin 
           xpc10 <= 10'd721/*721:xpc10:721*/;
           A_UINT[19'h6_1a80+10'h250] <= 32'd907627842;
           end 
          
      10'd721/*721:US*/:  begin 
           xpc10 <= 10'd722/*722:xpc10:722*/;
           A_UINT[19'h6_1a80+10'h254] <= 32'd853037301;
           end 
          
      10'd722/*722:US*/:  begin 
           xpc10 <= 10'd723/*723:xpc10:723*/;
           A_UINT[19'h6_1a80+10'h258] <= 32'd1067152940;
           end 
          
      10'd723/*723:US*/:  begin 
           xpc10 <= 10'd724/*724:xpc10:724*/;
           A_UINT[19'h6_1a80+10'h25c] <= 32'd995781531;
           end 
          
      10'd724/*724:US*/:  begin 
           xpc10 <= 10'd725/*725:xpc10:725*/;
           A_UINT[19'h6_1a80+10'h260] <= 32'd51762726;
           end 
          
      10'd725/*725:US*/:  begin 
           xpc10 <= 10'd726/*726:xpc10:726*/;
           A_UINT[19'h6_1a80+10'h264] <= 32'd131386257;
           end 
          
      10'd726/*726:US*/:  begin 
           xpc10 <= 10'd727/*727:xpc10:727*/;
           A_UINT[19'h6_1a80+10'h268] <= 32'd177728840;
           end 
          
      10'd727/*727:US*/:  begin 
           xpc10 <= 10'd728/*728:xpc10:728*/;
           A_UINT[19'h6_1a80+10'h26c] <= 32'd240578815;
           end 
          
      10'd728/*728:US*/:  begin 
           xpc10 <= 10'd729/*729:xpc10:729*/;
           A_UINT[19'h6_1a80+10'h270] <= 32'd269590778;
           end 
          
      10'd729/*729:US*/:  begin 
           xpc10 <= 10'd730/*730:xpc10:730*/;
           A_UINT[19'h6_1a80+10'h274] <= 32'd349224269;
           end 
          
      10'd730/*730:US*/:  begin 
           xpc10 <= 10'd731/*731:xpc10:731*/;
           A_UINT[19'h6_1a80+10'h278] <= 32'd429104020;
           end 
          
      10'd731/*731:US*/:  begin 
           xpc10 <= 10'd732/*732:xpc10:732*/;
           A_UINT[19'h6_1a80+10'h27c] <= 32'd491947555;
           end 
          
      10'd732/*732:US*/:  begin 
           xpc10 <= 10'd733/*733:xpc10:733*/;
           A_UINT[19'h6_1a80+10'h280] <= -32'd248556018;
           end 
          
      10'd733/*733:US*/:  begin 
           xpc10 <= 10'd734/*734:xpc10:734*/;
           A_UINT[19'h6_1a80+10'h284] <= -32'd168932423;
           end 
          
      10'd734/*734:US*/:  begin 
           xpc10 <= 10'd735/*735:xpc10:735*/;
           A_UINT[19'h6_1a80+10'h288] <= -32'd122852000;
           end 
          
      10'd735/*735:US*/:  begin 
           xpc10 <= 10'd736/*736:xpc10:736*/;
           A_UINT[19'h6_1a80+10'h28c] <= -32'd60002089;
           end 
          
      10'd736/*736:US*/:  begin 
           xpc10 <= 10'd737/*737:xpc10:737*/;
           A_UINT[19'h6_1a80+10'h290] <= -32'd500490030;
           end 
          
      10'd737/*737:US*/:  begin 
           xpc10 <= 10'd738/*738:xpc10:738*/;
           A_UINT[19'h6_1a80+10'h294] <= -32'd420856475;
           end 
          
      10'd738/*738:US*/:  begin 
           xpc10 <= 10'd739/*739:xpc10:739*/;
           A_UINT[19'h6_1a80+10'h298] <= -32'd341238852;
           end 
          
      10'd739/*739:US*/:  begin 
           xpc10 <= 10'd740/*740:xpc10:740*/;
           A_UINT[19'h6_1a80+10'h29c] <= -32'd278395381;
           end 
          
      10'd740/*740:US*/:  begin 
           xpc10 <= 10'd741/*741:xpc10:741*/;
           A_UINT[19'h6_1a80+10'h2a0] <= -32'd685261898;
           end 
          
      10'd741/*741:US*/:  begin 
           xpc10 <= 10'd742/*742:xpc10:742*/;
           A_UINT[19'h6_1a80+10'h2a4] <= -32'd739858943;
           end 
          
      10'd742/*742:US*/:  begin 
           xpc10 <= 10'd743/*743:xpc10:743*/;
           A_UINT[19'h6_1a80+10'h2a8] <= -32'd559578920;
           end 
          
      10'd743/*743:US*/:  begin 
           xpc10 <= 10'd744/*744:xpc10:744*/;
           A_UINT[19'h6_1a80+10'h2ac] <= -32'd630940305;
           end 
          
      10'd744/*744:US*/:  begin 
           xpc10 <= 10'd745/*745:xpc10:745*/;
           A_UINT[19'h6_1a80+10'h2b0] <= -32'd1004286614;
           end 
          
      10'd745/*745:US*/:  begin 
           xpc10 <= 10'd746/*746:xpc10:746*/;
           A_UINT[19'h6_1a80+10'h2b4] <= -32'd1058877219;
           end 
          
      10'd746/*746:US*/:  begin 
           xpc10 <= 10'd747/*747:xpc10:747*/;
           A_UINT[19'h6_1a80+10'h2b8] <= -32'd845023740;
           end 
          
      10'd747/*747:US*/:  begin 
           xpc10 <= 10'd748/*748:xpc10:748*/;
           A_UINT[19'h6_1a80+10'h2bc] <= -32'd916395085;
           end 
          
      10'd748/*748:US*/:  begin 
           xpc10 <= 10'd749/*749:xpc10:749*/;
           A_UINT[19'h6_1a80+10'h2c0] <= -32'd1119974018;
           end 
          
      10'd749/*749:US*/:  begin 
           xpc10 <= 10'd750/*750:xpc10:750*/;
           A_UINT[19'h6_1a80+10'h2c4] <= -32'd1174433591;
           end 
          
      10'd750/*750:US*/:  begin 
           xpc10 <= 10'd751/*751:xpc10:751*/;
           A_UINT[19'h6_1a80+10'h2c8] <= -32'd1262701040;
           end 
          
      10'd751/*751:US*/:  begin 
           xpc10 <= 10'd752/*752:xpc10:752*/;
           A_UINT[19'h6_1a80+10'h2cc] <= -32'd1333941337;
           end 
          
      10'd752/*752:US*/:  begin 
           xpc10 <= 10'd753/*753:xpc10:753*/;
           A_UINT[19'h6_1a80+10'h2d0] <= -32'd1371866206;
           end 
          
      10'd753/*753:US*/:  begin 
           xpc10 <= 10'd754/*754:xpc10:754*/;
           A_UINT[19'h6_1a80+10'h2d4] <= -32'd1426332139;
           end 
          
      10'd754/*754:US*/:  begin 
           xpc10 <= 10'd755/*755:xpc10:755*/;
           A_UINT[19'h6_1a80+10'h2d8] <= -32'd1481064244;
           end 
          
      10'd755/*755:US*/:  begin 
           xpc10 <= 10'd756/*756:xpc10:756*/;
           A_UINT[19'h6_1a80+10'h2dc] <= -32'd1552294533;
           end 
          
      10'd756/*756:US*/:  begin 
           xpc10 <= 10'd757/*757:xpc10:757*/;
           A_UINT[19'h6_1a80+10'h2e0] <= -32'd1690935098;
           end 
          
      10'd757/*757:US*/:  begin 
           xpc10 <= 10'd758/*758:xpc10:758*/;
           A_UINT[19'h6_1a80+10'h2e4] <= -32'd1611170447;
           end 
          
      10'd758/*758:US*/:  begin 
           xpc10 <= 10'd759/*759:xpc10:759*/;
           A_UINT[19'h6_1a80+10'h2e8] <= -32'd1833673816;
           end 
          
      10'd759/*759:US*/:  begin 
           xpc10 <= 10'd760/*760:xpc10:760*/;
           A_UINT[19'h6_1a80+10'h2ec] <= -32'd1770699233;
           end 
          
      10'd760/*760:US*/:  begin 
           xpc10 <= 10'd761/*761:xpc10:761*/;
           A_UINT[19'h6_1a80+10'h2f0] <= -32'd2009983462;
           end 
          
      10'd761/*761:US*/:  begin 
           xpc10 <= 10'd762/*762:xpc10:762*/;
           A_UINT[19'h6_1a80+10'h2f4] <= -32'd1930228819;
           end 
          
      10'd762/*762:US*/:  begin 
           xpc10 <= 10'd763/*763:xpc10:763*/;
           A_UINT[19'h6_1a80+10'h2f8] <= -32'd2119160460;
           end 
          
      10'd763/*763:US*/:  begin 
           xpc10 <= 10'd764/*764:xpc10:764*/;
           A_UINT[19'h6_1a80+10'h2fc] <= -32'd2056179517;
           end 
          
      10'd764/*764:US*/:  begin 
           xpc10 <= 10'd765/*765:xpc10:765*/;
           A_UINT[19'h6_1a80+10'h300] <= 32'd1569362073;
           end 
          
      10'd765/*765:US*/:  begin 
           xpc10 <= 10'd766/*766:xpc10:766*/;
           A_UINT[19'h6_1a80+10'h304] <= 32'd1498123566;
           end 
          
      10'd766/*766:US*/:  begin 
           xpc10 <= 10'd767/*767:xpc10:767*/;
           A_UINT[19'h6_1a80+10'h308] <= 32'd1409854455;
           end 
          
      10'd767/*767:US*/:  begin 
           xpc10 <= 10'd768/*768:xpc10:768*/;
           A_UINT[19'h6_1a80+10'h30c] <= 32'd1355396672;
           end 
          
      10'd768/*768:US*/:  begin 
           xpc10 <= 10'd769/*769:xpc10:769*/;
           A_UINT[19'h6_1a80+10'h310] <= 32'd1317987909;
           end 
          
      10'd769/*769:US*/:  begin 
           xpc10 <= 10'd770/*770:xpc10:770*/;
           A_UINT[19'h6_1a80+10'h314] <= 32'd1246755826;
           end 
          
      10'd770/*770:US*/:  begin 
           xpc10 <= 10'd771/*771:xpc10:771*/;
           A_UINT[19'h6_1a80+10'h318] <= 32'd1192025387;
           end 
          
      10'd771/*771:US*/:  begin 
           xpc10 <= 10'd772/*772:xpc10:772*/;
           A_UINT[19'h6_1a80+10'h31c] <= 32'd1137557660;
           end 
          
      10'd772/*772:US*/:  begin 
           xpc10 <= 10'd773/*773:xpc10:773*/;
           A_UINT[19'h6_1a80+10'h320] <= 32'd2072149281;
           end 
          
      10'd773/*773:US*/:  begin 
           xpc10 <= 10'd774/*774:xpc10:774*/;
           A_UINT[19'h6_1a80+10'h324] <= 32'd2135122070;
           end 
          
      10'd774/*774:US*/:  begin 
           xpc10 <= 10'd775/*775:xpc10:775*/;
           A_UINT[19'h6_1a80+10'h328] <= 32'd1912620623;
           end 
          
      10'd775/*775:US*/:  begin 
           xpc10 <= 10'd776/*776:xpc10:776*/;
           A_UINT[19'h6_1a80+10'h32c] <= 32'd1992383480;
           end 
          
      10'd776/*776:US*/:  begin 
           xpc10 <= 10'd777/*777:xpc10:777*/;
           A_UINT[19'h6_1a80+10'h330] <= 32'd1753615357;
           end 
          
      10'd777/*777:US*/:  begin 
           xpc10 <= 10'd778/*778:xpc10:778*/;
           A_UINT[19'h6_1a80+10'h334] <= 32'd1816598090;
           end 
          
      10'd778/*778:US*/:  begin 
           xpc10 <= 10'd779/*779:xpc10:779*/;
           A_UINT[19'h6_1a80+10'h338] <= 32'd1627664531;
           end 
          
      10'd779/*779:US*/:  begin 
           xpc10 <= 10'd780/*780:xpc10:780*/;
           A_UINT[19'h6_1a80+10'h33c] <= 32'd1707420964;
           end 
          
      10'd780/*780:US*/:  begin 
           xpc10 <= 10'd781/*781:xpc10:781*/;
           A_UINT[19'h6_1a80+10'h340] <= 32'd295390185;
           end 
          
      10'd781/*781:US*/:  begin 
           xpc10 <= 10'd782/*782:xpc10:782*/;
           A_UINT[19'h6_1a80+10'h344] <= 32'd358241886;
           end 
          
      10'd782/*782:US*/:  begin 
           xpc10 <= 10'd783/*783:xpc10:783*/;
           A_UINT[19'h6_1a80+10'h348] <= 32'd404320391;
           end 
          
      10'd783/*783:US*/:  begin 
           xpc10 <= 10'd784/*784:xpc10:784*/;
           A_UINT[19'h6_1a80+10'h34c] <= 32'd483945776;
           end 
          
      10'd784/*784:US*/:  begin 
           xpc10 <= 10'd785/*785:xpc10:785*/;
           A_UINT[19'h6_1a80+10'h350] <= 32'd43990325;
           end 
          
      10'd785/*785:US*/:  begin 
           xpc10 <= 10'd786/*786:xpc10:786*/;
           A_UINT[19'h6_1a80+10'h354] <= 32'd106832002;
           end 
          
      10'd786/*786:US*/:  begin 
           xpc10 <= 10'd787/*787:xpc10:787*/;
           A_UINT[19'h6_1a80+10'h358] <= 32'd186451547;
           end 
          
      10'd787/*787:US*/:  begin 
           xpc10 <= 10'd788/*788:xpc10:788*/;
           A_UINT[19'h6_1a80+10'h35c] <= 32'd266083308;
           end 
          
      10'd788/*788:US*/:  begin 
           xpc10 <= 10'd789/*789:xpc10:789*/;
           A_UINT[19'h6_1a80+10'h360] <= 32'd932423249;
           end 
          
      10'd789/*789:US*/:  begin 
           xpc10 <= 10'd790/*790:xpc10:790*/;
           A_UINT[19'h6_1a80+10'h364] <= 32'd861060070;
           end 
          
      10'd790/*790:US*/:  begin 
           xpc10 <= 10'd791/*791:xpc10:791*/;
           A_UINT[19'h6_1a80+10'h368] <= 32'd1041341759;
           end 
          
      10'd791/*791:US*/:  begin 
           xpc10 <= 10'd792/*792:xpc10:792*/;
           A_UINT[19'h6_1a80+10'h36c] <= 32'd986742920;
           end 
          
      10'd792/*792:US*/:  begin 
           xpc10 <= 10'd793/*793:xpc10:793*/;
           A_UINT[19'h6_1a80+10'h370] <= 32'd613929101;
           end 
          
      10'd793/*793:US*/:  begin 
           xpc10 <= 10'd794/*794:xpc10:794*/;
           A_UINT[19'h6_1a80+10'h374] <= 32'd542559546;
           end 
          
      10'd794/*794:US*/:  begin 
           xpc10 <= 10'd795/*795:xpc10:795*/;
           A_UINT[19'h6_1a80+10'h378] <= 32'd756411363;
           end 
          
      10'd795/*795:US*/:  begin 
           xpc10 <= 10'd796/*796:xpc10:796*/;
           A_UINT[19'h6_1a80+10'h37c] <= 32'd701822548;
           end 
          
      10'd796/*796:US*/:  begin 
           xpc10 <= 10'd797/*797:xpc10:797*/;
           A_UINT[19'h6_1a80+10'h380] <= -32'd978770311;
           end 
          
      10'd797/*797:US*/:  begin 
           xpc10 <= 10'd798/*798:xpc10:798*/;
           A_UINT[19'h6_1a80+10'h384] <= -32'd1050133554;
           end 
          
      10'd798/*798:US*/:  begin 
           xpc10 <= 10'd799/*799:xpc10:799*/;
           A_UINT[19'h6_1a80+10'h388] <= -32'd869589737;
           end 
          
      10'd799/*799:US*/:  begin 
           xpc10 <= 10'd800/*800:xpc10:800*/;
           A_UINT[19'h6_1a80+10'h38c] <= -32'd924188512;
           end 
          
      10'd800/*800:US*/:  begin 
           xpc10 <= 10'd801/*801:xpc10:801*/;
           A_UINT[19'h6_1a80+10'h390] <= -32'd693284699;
           end 
          
      10'd801/*801:US*/:  begin 
           xpc10 <= 10'd802/*802:xpc10:802*/;
           A_UINT[19'h6_1a80+10'h394] <= -32'd764654318;
           end 
          
      10'd802/*802:US*/:  begin 
           xpc10 <= 10'd803/*803:xpc10:803*/;
           A_UINT[19'h6_1a80+10'h398] <= -32'd550540341;
           end 
          
      10'd803/*803:US*/:  begin 
           xpc10 <= 10'd804/*804:xpc10:804*/;
           A_UINT[19'h6_1a80+10'h39c] <= -32'd605129092;
           end 
          
      10'd804/*804:US*/:  begin 
           xpc10 <= 10'd805/*805:xpc10:805*/;
           A_UINT[19'h6_1a80+10'h3a0] <= -32'd475935807;
           end 
          
      10'd805/*805:US*/:  begin 
           xpc10 <= 10'd806/*806:xpc10:806*/;
           A_UINT[19'h6_1a80+10'h3a4] <= -32'd413084042;
           end 
          
      10'd806/*806:US*/:  begin 
           xpc10 <= 10'd807/*807:xpc10:807*/;
           A_UINT[19'h6_1a80+10'h3a8] <= -32'd366743377;
           end 
          
      10'd807/*807:US*/:  begin 
           xpc10 <= 10'd808/*808:xpc10:808*/;
           A_UINT[19'h6_1a80+10'h3ac] <= -32'd287118056;
           end 
          
      10'd808/*808:US*/:  begin 
           xpc10 <= 10'd809/*809:xpc10:809*/;
           A_UINT[19'h6_1a80+10'h3b0] <= -32'd257573603;
           end 
          
      10'd809/*809:US*/:  begin 
           xpc10 <= 10'd810/*810:xpc10:810*/;
           A_UINT[19'h6_1a80+10'h3b4] <= -32'd194731862;
           end 
          
      10'd810/*810:US*/:  begin 
           xpc10 <= 10'd811/*811:xpc10:811*/;
           A_UINT[19'h6_1a80+10'h3b8] <= -32'd114850189;
           end 
          
      10'd811/*811:US*/:  begin 
           xpc10 <= 10'd812/*812:xpc10:812*/;
           A_UINT[19'h6_1a80+10'h3bc] <= -32'd35218492;
           end 
          
      10'd812/*812:US*/:  begin 
           xpc10 <= 10'd813/*813:xpc10:813*/;
           A_UINT[19'h6_1a80+10'h3c0] <= -32'd1984365303;
           end 
          
      10'd813/*813:US*/:  begin 
           xpc10 <= 10'd814/*814:xpc10:814*/;
           A_UINT[19'h6_1a80+10'h3c4] <= -32'd1921392450;
           end 
          
      10'd814/*814:US*/:  begin 
           xpc10 <= 10'd815/*815:xpc10:815*/;
           A_UINT[19'h6_1a80+10'h3c8] <= -32'd2143631769;
           end 
          
      10'd815/*815:US*/:  begin 
           xpc10 <= 10'd816/*816:xpc10:816*/;
           A_UINT[19'h6_1a80+10'h3cc] <= -32'd2063868976;
           end 
          
      10'd816/*816:US*/:  begin 
           xpc10 <= 10'd817/*817:xpc10:817*/;
           A_UINT[19'h6_1a80+10'h3d0] <= -32'd1698919467;
           end 
          
      10'd817/*817:US*/:  begin 
           xpc10 <= 10'd818/*818:xpc10:818*/;
           A_UINT[19'h6_1a80+10'h3d4] <= -32'd1635936670;
           end 
          
      10'd818/*818:US*/:  begin 
           xpc10 <= 10'd819/*819:xpc10:819*/;
           A_UINT[19'h6_1a80+10'h3d8] <= -32'd1824608069;
           end 
          
      10'd819/*819:US*/:  begin 
           xpc10 <= 10'd820/*820:xpc10:820*/;
           A_UINT[19'h6_1a80+10'h3dc] <= -32'd1744851700;
           end 
          
      10'd820/*820:US*/:  begin 
           xpc10 <= 10'd821/*821:xpc10:821*/;
           A_UINT[19'h6_1a80+10'h3e0] <= -32'd1347415887;
           end 
          
      10'd821/*821:US*/:  begin 
           xpc10 <= 10'd822/*822:xpc10:822*/;
           A_UINT[19'h6_1a80+10'h3e4] <= -32'd1418654458;
           end 
          
      10'd822/*822:US*/:  begin 
           xpc10 <= 10'd823/*823:xpc10:823*/;
           A_UINT[19'h6_1a80+10'h3e8] <= -32'd1506661409;
           end 
          
      10'd823/*823:US*/:  begin 
           xpc10 <= 10'd824/*824:xpc10:824*/;
           A_UINT[19'h6_1a80+10'h3ec] <= -32'd1561119128;
           end 
          
      10'd824/*824:US*/:  begin 
           xpc10 <= 10'd825/*825:xpc10:825*/;
           A_UINT[19'h6_1a80+10'h3f0] <= -32'd1129027987;
           end 
          
      10'd825/*825:US*/:  begin 
           xpc10 <= 10'd826/*826:xpc10:826*/;
           A_UINT[19'h6_1a80+10'h3f4] <= -32'd1200260134;
           end 
          
      10'd826/*826:US*/:  begin 
           xpc10 <= 10'd827/*827:xpc10:827*/;
           A_UINT[19'h6_1a80+10'h3f8] <= -32'd1254728445;
           end 
          
      10'd827/*827:US*/:  begin 
           xpc10 <= 10'd828/*828:xpc10:828*/;
           A_SINT[19'h6_266c+3'd4] <= 32'd78;
           A_UINT[19'h6_1a80+10'h3fc] <= -32'd1309196108;
           end 
          
      10'd828/*828:US*/:  begin 
           xpc10 <= 10'd829/*829:xpc10:829*/;
           A_SINT[19'h6_266c+4'd8] <= 32'd2;
           end 
          
      10'd829/*829:US*/:  begin 
           xpc10 <= 10'd830/*830:xpc10:830*/;
           A_SINT[19'h6_2b5c+3'd4] <= 32'd78;
           end 
          
      10'd830/*830:US*/:  begin 
           xpc10 <= 10'd831/*831:xpc10:831*/;
           A_SINT[19'h6_2b5c+4'd8] <= 32'd2;
           end 
          
      10'd831/*831:US*/:  begin 
           xpc10 <= 10'd832/*832:xpc10:832*/;
           A_SINT[19'h6_304c+3'd4] <= 32'd78;
           end 
          
      10'd832/*832:US*/:  begin 
           xpc10 <= 10'd833/*833:xpc10:833*/;
           A_SINT[19'h6_304c+4'd8] <= 32'd2;
           end 
          
      10'd833/*833:US*/:  begin 
           xpc10 <= 10'd834/*834:xpc10:834*/;
           A_SINT[19'h6_353c+3'd4] <= 32'd78;
           end 
          
      10'd839/*839:US*/:  begin 
           xpc10 <= 10'd840/*840:xpc10:840*/;
           TSPsw1_2_V_0 <= 32'd0;
           end 
          
      10'd840/*840:US*/: if ((TSPsw1_2_V_0<2'd2))  xpc10 <= 10'd861/*861:xpc10:861*/;
           else  begin 
               xpc10 <= 10'd841/*841:xpc10:841*/;
               TSPsw1_2_V_1 <= 32'd1;
               end 
              
      10'd841/*841:US*/: if ((TSPsw1_2_V_1<7'd78))  xpc10 <= 10'd857/*857:xpc10:857*/;
           else  begin 
               xpc10 <= 10'd842/*842:xpc10:842*/;
               TSPru0_12_V_1 <= 32'd0;
               end 
              
      10'd843/*843:US*/: if ((TSPen0_17_V_0<5'd20))  xpc10 <= 10'd856/*856:xpc10:856*/;
           else  begin 
               xpc10 <= 10'd844/*844:xpc10:844*/;
               TSPe0_SPILL_256 <= 32'd0;
               end 
              
      10'd844/*844:US*/:  begin 
           xpc10 <= 10'd845/*845:xpc10:845*/;
           TSPne2_10_V_3 <= 32'd0;
           TSPne2_10_V_2 <= TSPe0_SPILL_256;
           end 
          
      10'd848/*848:US*/: if ((TSPte2_13_V_2<7'h4d))  xpc10 <= 10'd849/*849:xpc10:849*/;
           else  begin 
               xpc10 <= 10'd846/*846:xpc10:846*/;
               TSPte2_13_V_0 <= 32'd1+TSPte2_13_V_0;
               end 
              
      10'd853/*853:US*/: if ((TSPne2_10_V_6<A_64_SS[64'h6_305c+64'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPne2_10_V_0
      )+(64'h_ffff_ffff_ffff_ffff&TSPne2_10_V_3))]))  begin 
               xpc10 <= 10'd854/*854:xpc10:854*/;
               TSPne2_10_V_6 <= A_64_SS[64'h6_305c+64'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPne2_10_V_0)+(64'h_ffff_ffff_ffff_ffff
              &TSPne2_10_V_3))];

               end 
               else  xpc10 <= 10'd854/*854:xpc10:854*/;

      10'd855/*855:US*/:  begin 
           xpc10 <= 10'd845/*845:xpc10:845*/;
           TSPne2_10_V_3 <= 1'd1+TSPne2_10_V_3;
           A_64_SS[19'h6_354c+4'h8*(A_SINT[19'h6_353c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPne2_10_V_1)+(64'h_ffff_ffff_ffff_ffff&1'd1+TSPne2_10_V_3
          ))] <= -64'd10+A_64_SS[64'h6_305c+64'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPne2_10_V_1)+(64'h_ffff_ffff_ffff_ffff
          &1'd1+TSPne2_10_V_3))];

           end 
          
      10'd857/*857:US*/:  begin 
           xpc10 <= 10'd858/*858:xpc10:858*/;
           A_64_SS[19'h6_267c+4'h8*(64'h_ffff_ffff_ffff_ffff&TSPsw1_2_V_1)] <= 64'd0;
           end 
          
      10'd858/*858:US*/:  begin 
           xpc10 <= 10'd859/*859:xpc10:859*/;
           A_64_SS[19'h6_2b6c+4'h8*(64'h_ffff_ffff_ffff_ffff&TSPsw1_2_V_1)] <= 64'd0;
           end 
          
      10'd859/*859:US*/:  begin 
           xpc10 <= 10'd860/*860:xpc10:860*/;
           A_64_SS[19'h6_305c+4'h8*(64'h_ffff_ffff_ffff_ffff&TSPsw1_2_V_1)] <= 64'd0;
           end 
          
      10'd860/*860:US*/:  begin 
           xpc10 <= 10'd841/*841:xpc10:841*/;
           TSPsw1_2_V_1 <= 32'd1+TSPsw1_2_V_1;
           A_64_SS[19'h6_354c+4'h8*(64'h_ffff_ffff_ffff_ffff&TSPsw1_2_V_1)] <= -64'd10;
           end 
          
      10'd861/*861:US*/:  begin 
           xpc10 <= 10'd862/*862:xpc10:862*/;
           d_monitor <= TSPsw1_2_V_0;
           A_64_SS[19'h6_267c+4'h8*A_SINT[19'h6_266c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPsw1_2_V_0)] <= 64'd0;
           end 
          
      10'd862/*862:US*/:  begin 
           xpc10 <= 10'd863/*863:xpc10:863*/;
           A_64_SS[19'h6_2b6c+4'h8*A_SINT[19'h6_2b5c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPsw1_2_V_0)] <= 64'd0;
           end 
          
      10'd863/*863:US*/:  begin 
           xpc10 <= 10'd864/*864:xpc10:864*/;
           A_64_SS[19'h6_305c+4'h8*A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPsw1_2_V_0)] <= 64'd0;
           end 
          
      10'd864/*864:US*/:  begin 
           xpc10 <= 10'd840/*840:xpc10:840*/;
           TSPsw1_2_V_0 <= 32'd1+TSPsw1_2_V_0;
           A_64_SS[19'h6_354c+4'h8*A_SINT[19'h6_353c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPsw1_2_V_0)] <= -64'd10;
           end 
          
      10'd865/*865:US*/: if ((TSPen1_8_V_0<5'd20))  xpc10 <= 10'd835/*835:xpc10:835*/;
           else  begin 
               xpc10 <= 10'd837/*837:xpc10:837*/;
               TSPe1_SPILL_256 <= 32'd0;
               end 
              endcase
      if ((xpc10==10'd835/*835:US*/))  xpc10 <= 10'd836/*836:xpc10:836*/;
          //End structure HPR sw_test.exe


       end 
      

assign hprpin256610 = A_64_SS[19'h6_354c+4'h8*(A_SINT[19'h6_353c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPne2_10_V_0)+(64'h_ffff_ffff_ffff_ffff&1'd1+TSPne2_10_V_3
))];

assign hprpin258710 = -3'd2+A_64_SS[19'h6_2b6c+4'h8*(A_SINT[19'h6_2b5c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPne2_10_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPne2_10_V_3
))];

assign hprpin529710 = 32'h_ffff_ffff&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1
))];

assign hprpin534210 = 19'h6_1a80+19'h4*(19'd255&((-32'd1&((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255&(hprpin529710>>>5'd16)))? -32'd1&((19'h6_3b60+4'd8==19'h6_1a80
+3'h4*(8'd255&((-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0
)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8
], 8'd0})>>5'd24)))? -32'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff
&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT
[19'h6_3b60+4'd8], 8'd0}: A_UINT[32'h6_1a80+3'h4*(8'd255&((-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c
+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60
+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0})>>5'd24))])^((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255&(hprpin529710>>>4'd8)))? -32'd1
&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff
&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT[32'h6_1a80
+3'h4*(8'd255&(hprpin529710>>>4'd8))])^{-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff
&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT
[19'h6_3b60+4'd8], 8'd0}, 8'd0}: A_UINT[32'h6_1a80+3'h4*(8'd255&(hprpin529710>>>5'd16))])^((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255&
((-2'd1&((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255&((-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+
3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60
+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0})>>5'd24)))? -32'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c
+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60
+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT[32'h6_1a80+3'h4*(8'd255&((-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c
+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80
+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0})>>5'd24))])^((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255
&(hprpin529710>>>4'd8)))? -32'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff
&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT
[19'h6_3b60+4'd8], 8'd0}: A_UINT[32'h6_1a80+3'h4*(8'd255&(hprpin529710>>>4'd8))])^{-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c
+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80
+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0}, 8'd0})>>5'd24)))? -32'd1&((19'h6_3b60+4'd8==19'h6_1a80
+3'h4*(8'd255&((-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0
)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8
], 8'd0})>>5'd24)))? -32'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff
&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT
[19'h6_3b60+4'd8], 8'd0}: A_UINT[32'h6_1a80+3'h4*(8'd255&((-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c
+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60
+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0})>>5'd24))])^((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255&(hprpin529710>>>4'd8)))? -32'd1
&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff
&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT[32'h6_1a80
+3'h4*(8'd255&(hprpin529710>>>4'd8))])^{-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff
&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT
[19'h6_3b60+4'd8], 8'd0}, 8'd0}: A_UINT[32'h6_1a80+3'h4*(8'd255&((-2'd1&((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255&((-2'd1&A_UINT[19'h6_1a80
+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1
))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0})>>5'd24)))? -32'd1&A_UINT[19'h6_1a80
+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1
))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT[32'h6_1a80+3'h4*(8'd255
&((-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff
&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0})>>5'd24))])^((19'h6_3b60
+4'd8==19'h6_1a80+3'h4*(8'd255&(hprpin529710>>>4'd8)))? -32'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c
+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60
+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT[32'h6_1a80+3'h4*(8'd255&(hprpin529710>>>4'd8))])^{-2'd1&A_UINT[19'h6_1a80+3'h4
*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1
))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0}, 8'd0})>>5'd24))])^{-2'd1&((19'h6_3b60
+4'd8==19'h6_1a80+3'h4*(8'd255&((-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff
&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT
[19'h6_3b60+4'd8], 8'd0})>>5'd24)))? -32'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff
&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT
[19'h6_3b60+4'd8], 8'd0}: A_UINT[32'h6_1a80+3'h4*(8'd255&((-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c
+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60
+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0})>>5'd24))])^((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255&(hprpin529710>>>4'd8)))? -32'd1
&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff
&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT[32'h6_1a80
+3'h4*(8'd255&(hprpin529710>>>4'd8))])^{-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff
&TSPcr2_16_V_0)+(64'h_ffff_ffff_ffff_ffff&TSPcr2_16_V_1))])]^A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^{A_UINT
[19'h6_3b60+4'd8], 8'd0}, 8'd0}, 8'd0})>>5'd24));

assign hprpin536910 = 32'h_ffff_ffff&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2
))];

assign hprpin540610 = 19'h6_1a80+19'h4*(19'd255&((-32'd1&((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255&((-2'd1&((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255&((-2'd1
&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c
+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0})>>5'd24)))? -2'd1
&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c
+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT[19'h6_1a80
+3'h4*(8'd255&((-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c
+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60
+4'd8], 8'd0})>>5'd24))])^((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255&(hprpin536910>>>4'd8)))? -2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT
[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff
&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT[19'h6_1a80+3'h4*(8'd255&(hprpin536910
>>>4'd8))])^{-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c
+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60
+4'd8], 8'd0}, 8'd0})>>5'd24)))? -32'd1&((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255&((-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60
+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1
)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0})>>5'd24)))? -2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT
[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff
&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT[19'h6_1a80+3'h4*(8'd255&((-2'd1&
A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c
+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0})>>5'd24))]
)^((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255&(hprpin536910>>>4'd8)))? -2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>
5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff
&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT[19'h6_1a80+3'h4*(8'd255&(hprpin536910>>>4'd8))])^{-2'd1&A_UINT[19'h6_1a80
+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff
&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0}, 8'd0}: A_UINT[32'h6_1a80+3'h4*(8'd255&((-2'd1
&((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255&((-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80
+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2
))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0})>>5'd24)))? -2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80
+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2
))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT[19'h6_1a80+3'h4*(8'd255&((-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]
>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff
&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0})>>5'd24))])^((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255&(hprpin536910>>>4'd8)))? -2'd1
&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c
+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT[19'h6_1a80
+3'h4*(8'd255&(hprpin536910>>>4'd8))])^{-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4
*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2
))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0}, 8'd0})>>5'd24))])^((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255&(hprpin536910>>>5'd16)))? -32'd1&
((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255&((-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80
+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2
))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0})>>5'd24)))? -2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80
+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2
))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT[19'h6_1a80+3'h4*(8'd255&((-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]
>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff
&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0})>>5'd24))])^((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255&(hprpin536910>>>4'd8)))? -2'd1
&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c
+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT[19'h6_1a80
+3'h4*(8'd255&(hprpin536910>>>4'd8))])^{-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4
*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2
))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0}, 8'd0}: A_UINT[32'h6_1a80+3'h4*(8'd255&(hprpin536910>>>5'd16))])^{-2'd1&((19'h6_3b60+4'd8==19'h6_1a80
+3'h4*(8'd255&((-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c
+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60
+4'd8], 8'd0})>>5'd24)))? -2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS
[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT
[19'h6_3b60+4'd8], 8'd0}: A_UINT[19'h6_1a80+3'h4*(8'd255&((-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT
[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff
&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0})>>5'd24))])^((19'h6_3b60+4'd8==19'h6_1a80+3'h4*(8'd255&(hprpin536910>>>4'd8)))? -2'd1
&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c
+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0}: A_UINT[19'h6_1a80
+3'h4*(8'd255&(hprpin536910>>>4'd8))])^{-2'd1&A_UINT[19'h6_1a80+3'h4*(8'd255&(A_UINT[19'h6_3b60+4'd8]>>5'd24))]^A_UINT[19'h6_1a80+3'h4
*(8'd255&A_64_SS[19'h6_305c+4'h8*(A_SINT[19'h6_304c+3'd4]*(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_1)+(64'h_ffff_ffff_ffff_ffff&TSPte2_13_V_2
))])]^{A_UINT[19'h6_3b60+4'd8], 8'd0}, 8'd0}, 8'd0})>>5'd24));

//Total area 0
// 1 vectors of width 10
// 1 vectors of width 64
// 576 bits in scalar variables
// Total state bits in module = 650 bits.
// 230 continuously assigned (wire/non-state) bits 
// Total number of leaf cells = 0
endmodule

//  
// LCP delay estimations included: turn off with -vnl-lcp-delay-estimate=disable
// eof (HPR L/S Verilog)
