

// CBG Orangepath HPR L/S System

// Verilog output file generated at 21/01/2016 13:21:23
// Kiwi Scientific Acceleration (KiwiC .net/CIL/C# to Verilog/SystemC compiler): Version alpha 2.01: January-2016 Unix 3.19.8.100
//  /home/djg11/d320/hprls/kiwipro/kiwic/distro/lib/kiwic.exe -verilog-roundtrip=disable -report-each-step -kiwic-finish=enable -kiwic-kcode-dump=enable -kiwic-cil-dump=separately -gtrace-loglevel=0 -restructure2=disable sw_test.exe -vnl=sw_test_a1 -sim 100000 -vnl-rootmodname=DUT -vnl-resets=synchronous -diosim-tl=100
`timescale 1ns/10ps


module DUT(output [31:0] result, output reg signed [63:0] d_monitor, output reg [31:0] phase, input clk, input reset);
  integer TSPru0_12_V_0;
  integer TSPru0_12_V_1;
  integer TSPin0_6_V_0;
  integer TSPen1_8_V_0;
  integer TSPsw1_2_V_0;
  integer TSPsw1_2_V_1;
  integer TSPne2_10_V_0;
  integer TSPne2_10_V_1;
  integer TSPne2_10_V_2;
  integer TSPne2_10_V_3;
  integer TSPne2_10_V_4;
  reg signed [63:0] TSPne2_10_V_7;
  integer TSPen0_17_V_0;
  integer TSPte2_13_V_0;
  integer TSPte2_13_V_1;
  integer TSPte2_13_V_2;
  integer TSPcr2_16_V_0;
  integer TSPcr2_16_V_1;
  reg signed [63:0] TSPcr2_16_V_2;
  reg [7:0] TCpr0_13_V_0;
  reg [7:0] TCpr0_21_V_0;
  reg [7:0] TCpr0_29_V_0;
  reg [7:0] TCpr0_35_V_0;
  reg [7:0] TCpr0_40_V_0;
  reg [7:0] TCpr0_44_V_0;
  integer TSPe1_SPILL_256;
  integer TSPe0_SPILL_256;
  reg signed [63:0] A_64_SS_CC_SCALbx52_ARA0[155:0];
  reg signed [63:0] A_64_SS_CC_SCALbx54_ARB0[155:0];
  reg signed [63:0] A_64_SS_CC_SCALbx56_ARC0[155:0];
  reg signed [63:0] A_64_SS_CC_SCALbx58_ARD0[155:0];
  reg [31:0] A_UINT_CC_SCALbx34_ARA0[509:0];
  reg [31:0] A_UINT_CC_SCALbx36_crc_reg;
  reg [31:0] A_UINT_CC_SCALbx36_byteno;
  reg [31:0] A_UINT_CC_SCALbx38_crc_reg;
  reg signed [31:0] A_SINT_CC_SCALbx16_ARA0[797:0];
  reg signed [31:0] A_SINT_CC_SCALbx32_d2dim0;
  reg signed [31:0] A_SINT_CC_SCALbx44_d2dim0;
  reg signed [31:0] A_SINT_CC_SCALbx40_d2dim0;
  reg signed [31:0] A_SINT_CC_SCALbx46_d2dim0;
  reg signed [31:0] A_SINT_CC_SCALbx26_ARJ0[76:0];
  reg signed [31:0] A_SINT_CC_SCALbx42_d2dim0;
  reg signed [15:0] A_16_SS_CC_SCALbx10_ARA0[147:0];
  reg signed [15:0] A_16_SS_CC_SCALbx12_ARB0[37:0];
  reg signed [15:0] A_16_SS_CC_SCALbx14_ARC0[151:0];
  reg [5:0] xpc10;
 always   @(posedge clk )  begin 
      //Start structure HPR sw_test.exe
      if (reset)  begin 
               A_SINT_CC_SCALbx40_d2dim0 <= 32'd0;
               A_SINT_CC_SCALbx42_d2dim0 <= 32'd0;
               A_SINT_CC_SCALbx44_d2dim0 <= 32'd0;
               A_SINT_CC_SCALbx46_d2dim0 <= 32'd0;
               A_SINT_CC_SCALbx32_d2dim0 <= 32'd0;
               TSPen1_8_V_0 <= 32'd0;
               TSPin0_6_V_0 <= 32'd0;
               TCpr0_40_V_0 <= 8'd0;
               TCpr0_44_V_0 <= 8'd0;
               A_UINT_CC_SCALbx38_crc_reg <= 32'd0;
               TSPru0_12_V_0 <= 32'd0;
               TSPne2_10_V_1 <= 32'd0;
               TSPne2_10_V_0 <= 32'd0;
               TSPne2_10_V_2 <= 32'd0;
               phase <= 32'd0;
               TSPte2_13_V_1 <= 32'd0;
               TSPcr2_16_V_0 <= 32'd0;
               TSPru0_12_V_1 <= 32'd0;
               TCpr0_13_V_0 <= 8'd0;
               TSPcr2_16_V_2 <= 64'd0;
               TCpr0_21_V_0 <= 8'd0;
               TCpr0_29_V_0 <= 8'd0;
               A_UINT_CC_SCALbx36_byteno <= 32'd0;
               TCpr0_35_V_0 <= 8'd0;
               TSPcr2_16_V_1 <= 32'd0;
               A_UINT_CC_SCALbx36_crc_reg <= 32'd0;
               TSPte2_13_V_0 <= 32'd0;
               TSPte2_13_V_2 <= 32'd0;
               TSPne2_10_V_4 <= 32'd0;
               TSPne2_10_V_7 <= 64'd0;
               TSPne2_10_V_3 <= 32'd0;
               TSPe0_SPILL_256 <= 32'd0;
               TSPen0_17_V_0 <= 32'd0;
               TSPsw1_2_V_1 <= 32'd0;
               TSPsw1_2_V_0 <= 32'd0;
               d_monitor <= 64'd0;
               TSPe1_SPILL_256 <= 32'd0;
               xpc10 <= 6'd0;
               end 
               else  begin 
              if ((xpc10==0/*0:US*/))  begin 
                      $display("Smith Waterman Simple Test Start. Iterations=%d", 33'h1ffffffff&32'd1);
                      $display("waypoint %d %d", 2'd2, 0);
                       end 
                      if (((33'h1ffffffff&32'd1+TSPin0_6_V_0)>=(33'h1ffffffff&32'h4d)) && (xpc10==2'd3/*3:US*/)) $display("waypoint %d %d"
                  , 2'd3, 0);
                  if ((TSPru0_12_V_0>=(33'h1ffffffff&32'd1)) && (xpc10==3'd4/*4:US*/))  begin 
                      $display("waypoint %d %d", 4'd12, 0);
                      $display("CRC RESET");
                      $display("crc reg now:  reg=%h", 33'h1ffffffff&-32'd1);
                       end 
                      
              case (xpc10)

              3'd7/*7:US*/: $display("self test startup %d a ", A_UINT_CC_SCALbx34_ARA0[32'd255]);

              4'd8/*8:US*/: $display("self test startup %d b ", 9'h1ff&8'd255);

              4'd9/*9:US*/: $display("self test startup %d c ", A_UINT_CC_SCALbx34_ARA0[32'd255]);

              4'd15/*15:US*/:  begin 
                  $display("self test yields %d (should be 821105832)", A_UINT_CC_SCALbx38_crc_reg);
                  $display("Smith Waterman Simple Test End.");
                  $finish(0);
                   end 
                  endcase
              if ((TSPru0_12_V_1<2'd3) && (xpc10==5'd19/*19:US*/))  begin 
                      $display("waypoint %d %d", 3'd6, TSPru0_12_V_1);
                      $display("waypoint %d %d", 3'd4, 0);
                       end 
                      if ((TSPne2_10_V_3>=(33'h1ffffffff&32'h4d)) && (xpc10==5'd22/*22:US*/))  begin 
                      $display("waypoint %d %d", 4'd8, TSPru0_12_V_1);
                      $display("Scored h matrix %d", TSPru0_12_V_1);
                       end 
                      if ((TSPte2_13_V_0>=2'd2) && (xpc10==5'd23/*23:US*/))  begin 
                      $display("waypoint %d %d", 4'd10, TSPru0_12_V_1);
                      $display("CRC RESET");
                      $display("crc reg now:  reg=%h", 33'h1ffffffff&-32'd1);
                       end 
                      
              case (xpc10)

              0/*0:US*/:  begin 
                   xpc10 <= 1'd1/*1:xpc10:1*/;
                   TSPen1_8_V_0 <= 33'h1ffffffff&32'd0;
                   TSPin0_6_V_0 <= 33'h1ffffffff&32'd0;
                   phase <= 33'h1ffffffff&32'd2;
                   A_SINT_CC_SCALbx40_d2dim0 <= 33'h1ffffffff&32'd78;
                   A_SINT_CC_SCALbx42_d2dim0 <= 33'h1ffffffff&32'd78;
                   A_SINT_CC_SCALbx44_d2dim0 <= 33'h1ffffffff&32'd78;
                   A_SINT_CC_SCALbx46_d2dim0 <= 33'h1ffffffff&32'd78;
                   A_SINT_CC_SCALbx32_d2dim0 <= 33'h1ffffffff&32'd20;
                   A_UINT_CC_SCALbx34_ARA0[32'd255] <= 33'h1ffffffff&-32'd1309196108;
                   A_UINT_CC_SCALbx34_ARA0[8'd254] <= 33'h1ffffffff&-32'd1254728445;
                   A_UINT_CC_SCALbx34_ARA0[8'd253] <= 33'h1ffffffff&-32'd1200260134;
                   A_UINT_CC_SCALbx34_ARA0[8'd252] <= 33'h1ffffffff&-32'd1129027987;
                   A_UINT_CC_SCALbx34_ARA0[8'd251] <= 33'h1ffffffff&-32'd1561119128;
                   A_UINT_CC_SCALbx34_ARA0[8'd250] <= 33'h1ffffffff&-32'd1506661409;
                   A_UINT_CC_SCALbx34_ARA0[8'd249] <= 33'h1ffffffff&-32'd1418654458;
                   A_UINT_CC_SCALbx34_ARA0[8'd248] <= 33'h1ffffffff&-32'd1347415887;
                   A_UINT_CC_SCALbx34_ARA0[8'd247] <= 33'h1ffffffff&-32'd1744851700;
                   A_UINT_CC_SCALbx34_ARA0[8'd246] <= 33'h1ffffffff&-32'd1824608069;
                   A_UINT_CC_SCALbx34_ARA0[8'd245] <= 33'h1ffffffff&-32'd1635936670;
                   A_UINT_CC_SCALbx34_ARA0[8'd244] <= 33'h1ffffffff&-32'd1698919467;
                   A_UINT_CC_SCALbx34_ARA0[8'd243] <= 33'h1ffffffff&-32'd2063868976;
                   A_UINT_CC_SCALbx34_ARA0[8'd242] <= 33'h1ffffffff&-32'd2143631769;
                   A_UINT_CC_SCALbx34_ARA0[8'd241] <= 33'h1ffffffff&-32'd1921392450;
                   A_UINT_CC_SCALbx34_ARA0[8'd240] <= 33'h1ffffffff&-32'd1984365303;
                   A_UINT_CC_SCALbx34_ARA0[8'd239] <= 33'h1ffffffff&-32'd35218492;
                   A_UINT_CC_SCALbx34_ARA0[8'd238] <= 33'h1ffffffff&-32'd114850189;
                   A_UINT_CC_SCALbx34_ARA0[8'd237] <= 33'h1ffffffff&-32'd194731862;
                   A_UINT_CC_SCALbx34_ARA0[8'd236] <= 33'h1ffffffff&-32'd257573603;
                   A_UINT_CC_SCALbx34_ARA0[8'd235] <= 33'h1ffffffff&-32'd287118056;
                   A_UINT_CC_SCALbx34_ARA0[8'd234] <= 33'h1ffffffff&-32'd366743377;
                   A_UINT_CC_SCALbx34_ARA0[8'd233] <= 33'h1ffffffff&-32'd413084042;
                   A_UINT_CC_SCALbx34_ARA0[8'd232] <= 33'h1ffffffff&-32'd475935807;
                   A_UINT_CC_SCALbx34_ARA0[8'd231] <= 33'h1ffffffff&-32'd605129092;
                   A_UINT_CC_SCALbx34_ARA0[8'd230] <= 33'h1ffffffff&-32'd550540341;
                   A_UINT_CC_SCALbx34_ARA0[8'd229] <= 33'h1ffffffff&-32'd764654318;
                   A_UINT_CC_SCALbx34_ARA0[8'd228] <= 33'h1ffffffff&-32'd693284699;
                   A_UINT_CC_SCALbx34_ARA0[8'd227] <= 33'h1ffffffff&-32'd924188512;
                   A_UINT_CC_SCALbx34_ARA0[8'd226] <= 33'h1ffffffff&-32'd869589737;
                   A_UINT_CC_SCALbx34_ARA0[8'd225] <= 33'h1ffffffff&-32'd1050133554;
                   A_UINT_CC_SCALbx34_ARA0[8'd224] <= 33'h1ffffffff&-32'd978770311;
                   A_UINT_CC_SCALbx34_ARA0[8'd223] <= 33'h1ffffffff&32'd701822548;
                   A_UINT_CC_SCALbx34_ARA0[8'd222] <= 33'h1ffffffff&32'd756411363;
                   A_UINT_CC_SCALbx34_ARA0[8'd221] <= 33'h1ffffffff&32'd542559546;
                   A_UINT_CC_SCALbx34_ARA0[8'd220] <= 33'h1ffffffff&32'd613929101;
                   A_UINT_CC_SCALbx34_ARA0[8'd219] <= 33'h1ffffffff&32'd986742920;
                   A_UINT_CC_SCALbx34_ARA0[8'd218] <= 33'h1ffffffff&32'd1041341759;
                   A_UINT_CC_SCALbx34_ARA0[8'd217] <= 33'h1ffffffff&32'd861060070;
                   A_UINT_CC_SCALbx34_ARA0[8'd216] <= 33'h1ffffffff&32'd932423249;
                   A_UINT_CC_SCALbx34_ARA0[8'd215] <= 33'h1ffffffff&32'd266083308;
                   A_UINT_CC_SCALbx34_ARA0[8'd214] <= 33'h1ffffffff&32'd186451547;
                   A_UINT_CC_SCALbx34_ARA0[8'd213] <= 33'h1ffffffff&32'd106832002;
                   A_UINT_CC_SCALbx34_ARA0[8'd212] <= 33'h1ffffffff&32'd43990325;
                   A_UINT_CC_SCALbx34_ARA0[8'd211] <= 33'h1ffffffff&32'd483945776;
                   A_UINT_CC_SCALbx34_ARA0[8'd210] <= 33'h1ffffffff&32'd404320391;
                   A_UINT_CC_SCALbx34_ARA0[8'd209] <= 33'h1ffffffff&32'd358241886;
                   A_UINT_CC_SCALbx34_ARA0[8'd208] <= 33'h1ffffffff&32'd295390185;
                   A_UINT_CC_SCALbx34_ARA0[8'd207] <= 33'h1ffffffff&32'd1707420964;
                   A_UINT_CC_SCALbx34_ARA0[8'd206] <= 33'h1ffffffff&32'd1627664531;
                   A_UINT_CC_SCALbx34_ARA0[8'd205] <= 33'h1ffffffff&32'd1816598090;
                   A_UINT_CC_SCALbx34_ARA0[8'd204] <= 33'h1ffffffff&32'd1753615357;
                   A_UINT_CC_SCALbx34_ARA0[8'd203] <= 33'h1ffffffff&32'd1992383480;
                   A_UINT_CC_SCALbx34_ARA0[8'd202] <= 33'h1ffffffff&32'd1912620623;
                   A_UINT_CC_SCALbx34_ARA0[8'd201] <= 33'h1ffffffff&32'd2135122070;
                   A_UINT_CC_SCALbx34_ARA0[8'd200] <= 33'h1ffffffff&32'd2072149281;
                   A_UINT_CC_SCALbx34_ARA0[8'd199] <= 33'h1ffffffff&32'd1137557660;
                   A_UINT_CC_SCALbx34_ARA0[8'd198] <= 33'h1ffffffff&32'd1192025387;
                   A_UINT_CC_SCALbx34_ARA0[8'd197] <= 33'h1ffffffff&32'd1246755826;
                   A_UINT_CC_SCALbx34_ARA0[8'd196] <= 33'h1ffffffff&32'd1317987909;
                   A_UINT_CC_SCALbx34_ARA0[8'd195] <= 33'h1ffffffff&32'd1355396672;
                   A_UINT_CC_SCALbx34_ARA0[8'd194] <= 33'h1ffffffff&32'd1409854455;
                   A_UINT_CC_SCALbx34_ARA0[8'd193] <= 33'h1ffffffff&32'd1498123566;
                   A_UINT_CC_SCALbx34_ARA0[8'd192] <= 33'h1ffffffff&32'd1569362073;
                   A_UINT_CC_SCALbx34_ARA0[8'd191] <= 33'h1ffffffff&-32'd2056179517;
                   A_UINT_CC_SCALbx34_ARA0[8'd190] <= 33'h1ffffffff&-32'd2119160460;
                   A_UINT_CC_SCALbx34_ARA0[8'd189] <= 33'h1ffffffff&-32'd1930228819;
                   A_UINT_CC_SCALbx34_ARA0[8'd188] <= 33'h1ffffffff&-32'd2009983462;
                   A_UINT_CC_SCALbx34_ARA0[8'd187] <= 33'h1ffffffff&-32'd1770699233;
                   A_UINT_CC_SCALbx34_ARA0[8'd186] <= 33'h1ffffffff&-32'd1833673816;
                   A_UINT_CC_SCALbx34_ARA0[8'd185] <= 33'h1ffffffff&-32'd1611170447;
                   A_UINT_CC_SCALbx34_ARA0[8'd184] <= 33'h1ffffffff&-32'd1690935098;
                   A_UINT_CC_SCALbx34_ARA0[8'd183] <= 33'h1ffffffff&-32'd1552294533;
                   A_UINT_CC_SCALbx34_ARA0[8'd182] <= 33'h1ffffffff&-32'd1481064244;
                   A_UINT_CC_SCALbx34_ARA0[8'd181] <= 33'h1ffffffff&-32'd1426332139;
                   A_UINT_CC_SCALbx34_ARA0[8'd180] <= 33'h1ffffffff&-32'd1371866206;
                   A_UINT_CC_SCALbx34_ARA0[8'd179] <= 33'h1ffffffff&-32'd1333941337;
                   A_UINT_CC_SCALbx34_ARA0[8'd178] <= 33'h1ffffffff&-32'd1262701040;
                   A_UINT_CC_SCALbx34_ARA0[8'd177] <= 33'h1ffffffff&-32'd1174433591;
                   A_UINT_CC_SCALbx34_ARA0[8'd176] <= 33'h1ffffffff&-32'd1119974018;
                   A_UINT_CC_SCALbx34_ARA0[8'd175] <= 33'h1ffffffff&-32'd916395085;
                   A_UINT_CC_SCALbx34_ARA0[8'd174] <= 33'h1ffffffff&-32'd845023740;
                   A_UINT_CC_SCALbx34_ARA0[8'd173] <= 33'h1ffffffff&-32'd1058877219;
                   A_UINT_CC_SCALbx34_ARA0[8'd172] <= 33'h1ffffffff&-32'd1004286614;
                   A_UINT_CC_SCALbx34_ARA0[8'd171] <= 33'h1ffffffff&-32'd630940305;
                   A_UINT_CC_SCALbx34_ARA0[8'd170] <= 33'h1ffffffff&-32'd559578920;
                   A_UINT_CC_SCALbx34_ARA0[8'd169] <= 33'h1ffffffff&-32'd739858943;
                   A_UINT_CC_SCALbx34_ARA0[8'd168] <= 33'h1ffffffff&-32'd685261898;
                   A_UINT_CC_SCALbx34_ARA0[8'd167] <= 33'h1ffffffff&-32'd278395381;
                   A_UINT_CC_SCALbx34_ARA0[8'd166] <= 33'h1ffffffff&-32'd341238852;
                   A_UINT_CC_SCALbx34_ARA0[8'd165] <= 33'h1ffffffff&-32'd420856475;
                   A_UINT_CC_SCALbx34_ARA0[8'd164] <= 33'h1ffffffff&-32'd500490030;
                   A_UINT_CC_SCALbx34_ARA0[8'd163] <= 33'h1ffffffff&-32'd60002089;
                   A_UINT_CC_SCALbx34_ARA0[8'd162] <= 33'h1ffffffff&-32'd122852000;
                   A_UINT_CC_SCALbx34_ARA0[8'd161] <= 33'h1ffffffff&-32'd168932423;
                   A_UINT_CC_SCALbx34_ARA0[8'd160] <= 33'h1ffffffff&-32'd248556018;
                   A_UINT_CC_SCALbx34_ARA0[8'd159] <= 33'h1ffffffff&32'd491947555;
                   A_UINT_CC_SCALbx34_ARA0[8'd158] <= 33'h1ffffffff&32'd429104020;
                   A_UINT_CC_SCALbx34_ARA0[8'd157] <= 33'h1ffffffff&32'd349224269;
                   A_UINT_CC_SCALbx34_ARA0[8'd156] <= 33'h1ffffffff&32'd269590778;
                   A_UINT_CC_SCALbx34_ARA0[8'd155] <= 33'h1ffffffff&32'd240578815;
                   A_UINT_CC_SCALbx34_ARA0[8'd154] <= 33'h1ffffffff&32'd177728840;
                   A_UINT_CC_SCALbx34_ARA0[8'd153] <= 33'h1ffffffff&32'd131386257;
                   A_UINT_CC_SCALbx34_ARA0[8'd152] <= 33'h1ffffffff&32'd51762726;
                   A_UINT_CC_SCALbx34_ARA0[8'd151] <= 33'h1ffffffff&32'd995781531;
                   A_UINT_CC_SCALbx34_ARA0[8'd150] <= 33'h1ffffffff&32'd1067152940;
                   A_UINT_CC_SCALbx34_ARA0[8'd149] <= 33'h1ffffffff&32'd853037301;
                   A_UINT_CC_SCALbx34_ARA0[8'd148] <= 33'h1ffffffff&32'd907627842;
                   A_UINT_CC_SCALbx34_ARA0[8'd147] <= 33'h1ffffffff&32'd677256519;
                   A_UINT_CC_SCALbx34_ARA0[8'd146] <= 33'h1ffffffff&32'd748617968;
                   A_UINT_CC_SCALbx34_ARA0[8'd145] <= 33'h1ffffffff&32'd568075817;
                   A_UINT_CC_SCALbx34_ARA0[8'd144] <= 33'h1ffffffff&32'd622672798;
                   A_UINT_CC_SCALbx34_ARA0[8'd143] <= 33'h1ffffffff&32'd1363369299;
                   A_UINT_CC_SCALbx34_ARA0[8'd142] <= 33'h1ffffffff&32'd1434599652;
                   A_UINT_CC_SCALbx34_ARA0[8'd141] <= 33'h1ffffffff&32'd1489069629;
                   A_UINT_CC_SCALbx34_ARA0[8'd140] <= 33'h1ffffffff&32'd1543535498;
                   A_UINT_CC_SCALbx34_ARA0[8'd139] <= 33'h1ffffffff&32'd1111960463;
                   A_UINT_CC_SCALbx34_ARA0[8'd138] <= 33'h1ffffffff&32'd1183200824;
                   A_UINT_CC_SCALbx34_ARA0[8'd137] <= 33'h1ffffffff&32'd1271206113;
                   A_UINT_CC_SCALbx34_ARA0[8'd136] <= 33'h1ffffffff&32'd1325665622;
                   A_UINT_CC_SCALbx34_ARA0[8'd135] <= 33'h1ffffffff&32'd2001449195;
                   A_UINT_CC_SCALbx34_ARA0[8'd134] <= 33'h1ffffffff&32'd1938468188;
                   A_UINT_CC_SCALbx34_ARA0[8'd133] <= 33'h1ffffffff&32'd2127137669;
                   A_UINT_CC_SCALbx34_ARA0[8'd132] <= 33'h1ffffffff&32'd2047383090;
                   A_UINT_CC_SCALbx34_ARA0[8'd131] <= 33'h1ffffffff&32'd1682949687;
                   A_UINT_CC_SCALbx34_ARA0[8'd130] <= 33'h1ffffffff&32'd1619975040;
                   A_UINT_CC_SCALbx34_ARA0[8'd129] <= 33'h1ffffffff&32'd1842216281;
                   A_UINT_CC_SCALbx34_ARA0[32'd128] <= 33'h1ffffffff&32'd1762451694;
                   A_UINT_CC_SCALbx34_ARA0[7'd127] <= 33'h1ffffffff&-32'd654598054;
                   A_UINT_CC_SCALbx34_ARA0[7'd126] <= 33'h1ffffffff&-32'd600130067;
                   A_UINT_CC_SCALbx34_ARA0[7'd125] <= 33'h1ffffffff&-32'd780559564;
                   A_UINT_CC_SCALbx34_ARA0[7'd124] <= 33'h1ffffffff&-32'd709327229;
                   A_UINT_CC_SCALbx34_ARA0[7'd123] <= 33'h1ffffffff&-32'd872425850;
                   A_UINT_CC_SCALbx34_ARA0[7'd122] <= 33'h1ffffffff&-32'd817968335;
                   A_UINT_CC_SCALbx34_ARA0[7'd121] <= 33'h1ffffffff&-32'd1031934488;
                   A_UINT_CC_SCALbx34_ARA0[7'd120] <= 33'h1ffffffff&-32'd960696225;
                   A_UINT_CC_SCALbx34_ARA0[7'd119] <= 33'h1ffffffff&-32'd17609246;
                   A_UINT_CC_SCALbx34_ARA0[7'd118] <= 33'h1ffffffff&-32'd97365931;
                   A_UINT_CC_SCALbx34_ARA0[7'd117] <= 33'h1ffffffff&-32'd143559028;
                   A_UINT_CC_SCALbx34_ARA0[7'd116] <= 33'h1ffffffff&-32'd206542021;
                   A_UINT_CC_SCALbx34_ARA0[7'd115] <= 33'h1ffffffff&-32'd302564546;
                   A_UINT_CC_SCALbx34_ARA0[7'd114] <= 33'h1ffffffff&-32'd382327159;
                   A_UINT_CC_SCALbx34_ARA0[7'd113] <= 33'h1ffffffff&-32'd462094256;
                   A_UINT_CC_SCALbx34_ARA0[7'd112] <= 33'h1ffffffff&-32'd525066777;
                   A_UINT_CC_SCALbx34_ARA0[7'd111] <= 33'h1ffffffff&-32'd1796572374;
                   A_UINT_CC_SCALbx34_ARA0[7'd110] <= 33'h1ffffffff&-32'd1876203875;
                   A_UINT_CC_SCALbx34_ARA0[7'd109] <= 33'h1ffffffff&-32'd1654112188;
                   A_UINT_CC_SCALbx34_ARA0[7'd108] <= 33'h1ffffffff&-32'd1716953613;
                   A_UINT_CC_SCALbx34_ARA0[7'd107] <= 33'h1ffffffff&-32'd2014441994;
                   A_UINT_CC_SCALbx34_ARA0[7'd106] <= 33'h1ffffffff&-32'd2094067647;
                   A_UINT_CC_SCALbx34_ARA0[7'd105] <= 33'h1ffffffff&-32'd1905510760;
                   A_UINT_CC_SCALbx34_ARA0[7'd104] <= 33'h1ffffffff&-32'd1968362705;
                   A_UINT_CC_SCALbx34_ARA0[7'd103] <= 33'h1ffffffff&-32'd1293773166;
                   A_UINT_CC_SCALbx34_ARA0[7'd102] <= 33'h1ffffffff&-32'd1239184603;
                   A_UINT_CC_SCALbx34_ARA0[7'd101] <= 33'h1ffffffff&-32'd1151291908;
                   A_UINT_CC_SCALbx34_ARA0[7'd100] <= 33'h1ffffffff&-32'd1079922613;
                   A_UINT_CC_SCALbx34_ARA0[7'd99] <= 33'h1ffffffff&-32'd1578704818;
                   A_UINT_CC_SCALbx34_ARA0[7'd98] <= 33'h1ffffffff&-32'd1524105735;
                   A_UINT_CC_SCALbx34_ARA0[7'd97] <= 33'h1ffffffff&-32'd1469785312;
                   A_UINT_CC_SCALbx34_ARA0[7'd96] <= 33'h1ffffffff&-32'd1398421865;
                   A_UINT_CC_SCALbx34_ARA0[7'd95] <= 33'h1ffffffff&32'd1087903418;
                   A_UINT_CC_SCALbx34_ARA0[7'd94] <= 33'h1ffffffff&32'd1142491917;
                   A_UINT_CC_SCALbx34_ARA0[7'd93] <= 33'h1ffffffff&32'd1230646740;
                   A_UINT_CC_SCALbx34_ARA0[7'd92] <= 33'h1ffffffff&32'd1302016099;
                   A_UINT_CC_SCALbx34_ARA0[7'd91] <= 33'h1ffffffff&32'd1406951526;
                   A_UINT_CC_SCALbx34_ARA0[7'd90] <= 33'h1ffffffff&32'd1461550545;
                   A_UINT_CC_SCALbx34_ARA0[7'd89] <= 33'h1ffffffff&32'd1516133128;
                   A_UINT_CC_SCALbx34_ARA0[7'd88] <= 33'h1ffffffff&32'd1587496639;
                   A_UINT_CC_SCALbx34_ARA0[7'd87] <= 33'h1ffffffff&32'd1724971778;
                   A_UINT_CC_SCALbx34_ARA0[7'd86] <= 33'h1ffffffff&32'd1645340341;
                   A_UINT_CC_SCALbx34_ARA0[7'd85] <= 33'h1ffffffff&32'd1867694188;
                   A_UINT_CC_SCALbx34_ARA0[7'd84] <= 33'h1ffffffff&32'd1804852699;
                   A_UINT_CC_SCALbx34_ARA0[7'd83] <= 33'h1ffffffff&32'd1976864222;
                   A_UINT_CC_SCALbx34_ARA0[7'd82] <= 33'h1ffffffff&32'd1897238633;
                   A_UINT_CC_SCALbx34_ARA0[7'd81] <= 33'h1ffffffff&32'd2086057648;
                   A_UINT_CC_SCALbx34_ARA0[7'd80] <= 33'h1ffffffff&32'd2023205639;
                   A_UINT_CC_SCALbx34_ARA0[7'd79] <= 33'h1ffffffff&32'd214552010;
                   A_UINT_CC_SCALbx34_ARA0[7'd78] <= 33'h1ffffffff&32'd134795389;
                   A_UINT_CC_SCALbx34_ARA0[7'd77] <= 33'h1ffffffff&32'd88864420;
                   A_UINT_CC_SCALbx34_ARA0[7'd76] <= 33'h1ffffffff&32'd25881363;
                   A_UINT_CC_SCALbx34_ARA0[7'd75] <= 33'h1ffffffff&32'd533576470;
                   A_UINT_CC_SCALbx34_ARA0[7'd74] <= 33'h1ffffffff&32'd453813921;
                   A_UINT_CC_SCALbx34_ARA0[7'd73] <= 33'h1ffffffff&32'd374308984;
                   A_UINT_CC_SCALbx34_ARA0[7'd72] <= 33'h1ffffffff&32'd311336399;
                   A_UINT_CC_SCALbx34_ARA0[7'd71] <= 33'h1ffffffff&32'd717299826;
                   A_UINT_CC_SCALbx34_ARA0[7'd70] <= 33'h1ffffffff&32'd771767749;
                   A_UINT_CC_SCALbx34_ARA0[7'd69] <= 33'h1ffffffff&32'd591600412;
                   A_UINT_CC_SCALbx34_ARA0[7'd68] <= 33'h1ffffffff&32'd662832811;
                   A_UINT_CC_SCALbx34_ARA0[7'd67] <= 33'h1ffffffff&32'd969234094;
                   A_UINT_CC_SCALbx34_ARA0[7'd66] <= 33'h1ffffffff&32'd1023691545;
                   A_UINT_CC_SCALbx34_ARA0[7'd65] <= 33'h1ffffffff&32'd809987520;
                   A_UINT_CC_SCALbx34_ARA0[7'd64] <= 33'h1ffffffff&32'd881225847;
                   A_UINT_CC_SCALbx34_ARA0[6'd63] <= 33'h1ffffffff&-32'd327299027;
                   A_UINT_CC_SCALbx34_ARA0[6'd62] <= 33'h1ffffffff&-32'd390279782;
                   A_UINT_CC_SCALbx34_ARA0[6'd61] <= 33'h1ffffffff&-32'd436212925;
                   A_UINT_CC_SCALbx34_ARA0[6'd60] <= 33'h1ffffffff&-32'd515967244;
                   A_UINT_CC_SCALbx34_ARA0[6'd59] <= 33'h1ffffffff&-32'd8804623;
                   A_UINT_CC_SCALbx34_ARA0[6'd58] <= 33'h1ffffffff&-32'd71779514;
                   A_UINT_CC_SCALbx34_ARA0[6'd57] <= 33'h1ffffffff&-32'd151282273;
                   A_UINT_CC_SCALbx34_ARA0[6'd56] <= 33'h1ffffffff&-32'd231047128;
                   A_UINT_CC_SCALbx34_ARA0[6'd55] <= 33'h1ffffffff&-32'd898286187;
                   A_UINT_CC_SCALbx34_ARA0[6'd54] <= 33'h1ffffffff&-32'd827056094;
                   A_UINT_CC_SCALbx34_ARA0[6'd53] <= 33'h1ffffffff&-32'd1007220997;
                   A_UINT_CC_SCALbx34_ARA0[6'd52] <= 33'h1ffffffff&-32'd952755380;
                   A_UINT_CC_SCALbx34_ARA0[6'd51] <= 33'h1ffffffff&-32'd646886583;
                   A_UINT_CC_SCALbx34_ARA0[6'd50] <= 33'h1ffffffff&-32'd575645954;
                   A_UINT_CC_SCALbx34_ARA0[6'd49] <= 33'h1ffffffff&-32'd789352409;
                   A_UINT_CC_SCALbx34_ARA0[6'd48] <= 33'h1ffffffff&-32'd734892656;
                   A_UINT_CC_SCALbx34_ARA0[6'd47] <= 33'h1ffffffff&-32'd1603531939;
                   A_UINT_CC_SCALbx34_ARA0[6'd46] <= 33'h1ffffffff&-32'd1532160278;
                   A_UINT_CC_SCALbx34_ARA0[6'd45] <= 33'h1ffffffff&-32'd1444007885;
                   A_UINT_CC_SCALbx34_ARA0[6'd44] <= 33'h1ffffffff&-32'd1389417084;
                   A_UINT_CC_SCALbx34_ARA0[6'd43] <= 33'h1ffffffff&-32'd1284997759;
                   A_UINT_CC_SCALbx34_ARA0[6'd42] <= 33'h1ffffffff&-32'd1213636554;
                   A_UINT_CC_SCALbx34_ARA0[6'd41] <= 33'h1ffffffff&-32'd1159051537;
                   A_UINT_CC_SCALbx34_ARA0[6'd40] <= 33'h1ffffffff&-32'd1104454824;
                   A_UINT_CC_SCALbx34_ARA0[6'd39] <= 33'h1ffffffff&-32'd2040207643;
                   A_UINT_CC_SCALbx34_ARA0[6'd38] <= 33'h1ffffffff&-32'd2103051438;
                   A_UINT_CC_SCALbx34_ARA0[6'd37] <= 33'h1ffffffff&-32'd1880695413;
                   A_UINT_CC_SCALbx34_ARA0[6'd36] <= 33'h1ffffffff&-32'd1960329156;
                   A_UINT_CC_SCALbx34_ARA0[6'd35] <= 33'h1ffffffff&-32'd1788833735;
                   A_UINT_CC_SCALbx34_ARA0[6'd34] <= 33'h1ffffffff&-32'd1851683442;
                   A_UINT_CC_SCALbx34_ARA0[6'd33] <= 33'h1ffffffff&-32'd1662866601;
                   A_UINT_CC_SCALbx34_ARA0[6'd32] <= 33'h1ffffffff&-32'd1742489888;
                   A_UINT_CC_SCALbx34_ARA0[5'd31] <= 33'h1ffffffff&32'd1952343757;
                   A_UINT_CC_SCALbx34_ARA0[5'd30] <= 33'h1ffffffff&32'd1889500026;
                   A_UINT_CC_SCALbx34_ARA0[5'd29] <= 33'h1ffffffff&32'd2111593891;
                   A_UINT_CC_SCALbx34_ARA0[5'd28] <= 33'h1ffffffff&32'd2031960084;
                   A_UINT_CC_SCALbx34_ARA0[5'd27] <= 33'h1ffffffff&32'd1733955601;
                   A_UINT_CC_SCALbx34_ARA0[5'd26] <= 33'h1ffffffff&32'd1671105958;
                   A_UINT_CC_SCALbx34_ARA0[5'd25] <= 33'h1ffffffff&32'd1859660671;
                   A_UINT_CC_SCALbx34_ARA0[5'd24] <= 33'h1ffffffff&32'd1780037320;
                   A_UINT_CC_SCALbx34_ARA0[5'd23] <= 33'h1ffffffff&32'd1381403509;
                   A_UINT_CC_SCALbx34_ARA0[5'd22] <= 33'h1ffffffff&32'd1452775106;
                   A_UINT_CC_SCALbx34_ARA0[5'd21] <= 33'h1ffffffff&32'd1540665371;
                   A_UINT_CC_SCALbx34_ARA0[5'd20] <= 33'h1ffffffff&32'd1595256236;
                   A_UINT_CC_SCALbx34_ARA0[5'd19] <= 33'h1ffffffff&32'd1095957929;
                   A_UINT_CC_SCALbx34_ARA0[5'd18] <= 33'h1ffffffff&32'd1167319070;
                   A_UINT_CC_SCALbx34_ARA0[5'd17] <= 33'h1ffffffff&32'd1221641927;
                   A_UINT_CC_SCALbx34_ARA0[5'd16] <= 33'h1ffffffff&32'd1276238704;
                   A_UINT_CC_SCALbx34_ARA0[4'd15] <= 33'h1ffffffff&32'd944750013;
                   A_UINT_CC_SCALbx34_ARA0[4'd14] <= 33'h1ffffffff&32'd1015980042;
                   A_UINT_CC_SCALbx34_ARA0[4'd13] <= 33'h1ffffffff&32'd835552979;
                   A_UINT_CC_SCALbx34_ARA0[4'd12] <= 33'h1ffffffff&32'd890018660;
                   A_UINT_CC_SCALbx34_ARA0[4'd11] <= 33'h1ffffffff&32'd726387553;
                   A_UINT_CC_SCALbx34_ARA0[4'd10] <= 33'h1ffffffff&32'd797628118;
                   A_UINT_CC_SCALbx34_ARA0[4'd9] <= 33'h1ffffffff&32'd583659535;
                   A_UINT_CC_SCALbx34_ARA0[4'd8] <= 33'h1ffffffff&32'd638119352;
                   A_UINT_CC_SCALbx34_ARA0[3'd7] <= 33'h1ffffffff&32'd507990021;
                   A_UINT_CC_SCALbx34_ARA0[3'd6] <= 33'h1ffffffff&32'd445009330;
                   A_UINT_CC_SCALbx34_ARA0[3'd5] <= 33'h1ffffffff&32'd398814059;
                   A_UINT_CC_SCALbx34_ARA0[3'd4] <= 33'h1ffffffff&32'd319059676;
                   A_UINT_CC_SCALbx34_ARA0[2'd3] <= 33'h1ffffffff&32'd222504665;
                   A_UINT_CC_SCALbx34_ARA0[2'd2] <= 33'h1ffffffff&32'd159529838;
                   A_UINT_CC_SCALbx34_ARA0[32'd1] <= 33'h1ffffffff&32'd79764919;
                   A_UINT_CC_SCALbx34_ARA0[0] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[9'd399] <= 33'h1ffffffff&32'd10;
                   A_SINT_CC_SCALbx16_ARA0[9'd398] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[9'd397] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[9'd396] <= 33'h1ffffffff&-32'd3;
                   A_SINT_CC_SCALbx16_ARA0[9'd395] <= 33'h1ffffffff&-32'd3;
                   A_SINT_CC_SCALbx16_ARA0[9'd394] <= 33'h1ffffffff&-32'd4;
                   A_SINT_CC_SCALbx16_ARA0[9'd393] <= 33'h1ffffffff&-32'd4;
                   A_SINT_CC_SCALbx16_ARA0[9'd392] <= 33'h1ffffffff&-32'd5;
                   A_SINT_CC_SCALbx16_ARA0[9'd391] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[9'd390] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[9'd389] <= 33'h1ffffffff&-32'd1;
                   A_SINT_CC_SCALbx16_ARA0[9'd388] <= 33'h1ffffffff&-32'd4;
                   A_SINT_CC_SCALbx16_ARA0[9'd387] <= 33'h1ffffffff&-32'd1;
                   A_SINT_CC_SCALbx16_ARA0[9'd386] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[9'd385] <= 33'h1ffffffff&-32'd5;
                   A_SINT_CC_SCALbx16_ARA0[9'd384] <= 33'h1ffffffff&32'd7;
                   A_SINT_CC_SCALbx16_ARA0[9'd383] <= 33'h1ffffffff&-32'd4;
                   A_SINT_CC_SCALbx16_ARA0[9'd382] <= 33'h1ffffffff&-32'd4;
                   A_SINT_CC_SCALbx16_ARA0[9'd381] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[9'd380] <= 33'h1ffffffff&-32'd3;
                   A_SINT_CC_SCALbx16_ARA0[9'd379] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[9'd378] <= 33'h1ffffffff&32'd17;
                   A_SINT_CC_SCALbx16_ARA0[9'd377] <= 33'h1ffffffff&-32'd6;
                   A_SINT_CC_SCALbx16_ARA0[9'd376] <= 33'h1ffffffff&-32'd5;
                   A_SINT_CC_SCALbx16_ARA0[9'd375] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[9'd374] <= 33'h1ffffffff&32'd2;
                   A_SINT_CC_SCALbx16_ARA0[9'd373] <= 33'h1ffffffff&-32'd5;
                   A_SINT_CC_SCALbx16_ARA0[9'd372] <= 33'h1ffffffff&-32'd6;
                   A_SINT_CC_SCALbx16_ARA0[9'd371] <= 33'h1ffffffff&-32'd4;
                   A_SINT_CC_SCALbx16_ARA0[9'd370] <= 33'h1ffffffff&-32'd4;
                   A_SINT_CC_SCALbx16_ARA0[9'd369] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[9'd368] <= 33'h1ffffffff&-32'd3;
                   A_SINT_CC_SCALbx16_ARA0[9'd367] <= 33'h1ffffffff&-32'd5;
                   A_SINT_CC_SCALbx16_ARA0[9'd366] <= 33'h1ffffffff&-32'd3;
                   A_SINT_CC_SCALbx16_ARA0[9'd365] <= 33'h1ffffffff&-32'd7;
                   A_SINT_CC_SCALbx16_ARA0[9'd364] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[9'd363] <= 33'h1ffffffff&-32'd7;
                   A_SINT_CC_SCALbx16_ARA0[9'd362] <= 33'h1ffffffff&-32'd7;
                   A_SINT_CC_SCALbx16_ARA0[9'd361] <= 33'h1ffffffff&-32'd8;
                   A_SINT_CC_SCALbx16_ARA0[9'd360] <= 33'h1ffffffff&-32'd6;
                   A_SINT_CC_SCALbx16_ARA0[9'd359] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[9'd358] <= 33'h1ffffffff&-32'd6;
                   A_SINT_CC_SCALbx16_ARA0[9'd357] <= 33'h1ffffffff&32'd4;
                   A_SINT_CC_SCALbx16_ARA0[9'd356] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[9'd355] <= 33'h1ffffffff&-32'd1;
                   A_SINT_CC_SCALbx16_ARA0[9'd354] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[9'd353] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[9'd352] <= 33'h1ffffffff&-32'd1;
                   A_SINT_CC_SCALbx16_ARA0[9'd351] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[9'd350] <= 33'h1ffffffff&32'd2;
                   A_SINT_CC_SCALbx16_ARA0[9'd349] <= 33'h1ffffffff&32'd2;
                   A_SINT_CC_SCALbx16_ARA0[9'd348] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[9'd347] <= 33'h1ffffffff&32'd4;
                   A_SINT_CC_SCALbx16_ARA0[9'd346] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[9'd345] <= 33'h1ffffffff&-32'd1;
                   A_SINT_CC_SCALbx16_ARA0[9'd344] <= 33'h1ffffffff&-32'd1;
                   A_SINT_CC_SCALbx16_ARA0[9'd343] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[9'd342] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[9'd341] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[9'd340] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[9'd339] <= 33'h1ffffffff&-32'd3;
                   A_SINT_CC_SCALbx16_ARA0[9'd338] <= 33'h1ffffffff&-32'd5;
                   A_SINT_CC_SCALbx16_ARA0[9'd337] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[9'd336] <= 33'h1ffffffff&32'd3;
                   A_SINT_CC_SCALbx16_ARA0[9'd335] <= 33'h1ffffffff&32'd1;
                   A_SINT_CC_SCALbx16_ARA0[9'd334] <= 33'h1ffffffff&-32'd1;
                   A_SINT_CC_SCALbx16_ARA0[9'd333] <= 33'h1ffffffff&-32'd1;
                   A_SINT_CC_SCALbx16_ARA0[9'd332] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[9'd331] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[9'd330] <= 33'h1ffffffff&-32'd1;
                   A_SINT_CC_SCALbx16_ARA0[9'd329] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[9'd328] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[9'd327] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[9'd326] <= 33'h1ffffffff&-32'd1;
                   A_SINT_CC_SCALbx16_ARA0[9'd325] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[9'd324] <= 33'h1ffffffff&-32'd3;
                   A_SINT_CC_SCALbx16_ARA0[9'd323] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[9'd322] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[9'd321] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[9'd320] <= 33'h1ffffffff&32'd1;
                   A_SINT_CC_SCALbx16_ARA0[9'd319] <= 33'h1ffffffff&-32'd3;
                   A_SINT_CC_SCALbx16_ARA0[9'd318] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[9'd317] <= 33'h1ffffffff&-32'd1;
                   A_SINT_CC_SCALbx16_ARA0[9'd316] <= 33'h1ffffffff&32'd1;
                   A_SINT_CC_SCALbx16_ARA0[9'd315] <= 33'h1ffffffff&32'd2;
                   A_SINT_CC_SCALbx16_ARA0[9'd314] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[9'd313] <= 33'h1ffffffff&-32'd1;
                   A_SINT_CC_SCALbx16_ARA0[9'd312] <= 33'h1ffffffff&32'd1;
                   A_SINT_CC_SCALbx16_ARA0[9'd311] <= 33'h1ffffffff&32'd1;
                   A_SINT_CC_SCALbx16_ARA0[9'd310] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[9'd309] <= 33'h1ffffffff&-32'd3;
                   A_SINT_CC_SCALbx16_ARA0[9'd308] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[9'd307] <= 33'h1ffffffff&-32'd1;
                   A_SINT_CC_SCALbx16_ARA0[9'd306] <= 33'h1ffffffff&-32'd1;
                   A_SINT_CC_SCALbx16_ARA0[9'd305] <= 33'h1ffffffff&32'd1;
                   A_SINT_CC_SCALbx16_ARA0[9'd304] <= 33'h1ffffffff&-32'd3;
                   A_SINT_CC_SCALbx16_ARA0[9'd303] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[9'd302] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[9'd301] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[9'd300] <= 33'h1ffffffff&32'd1;
                   A_SINT_CC_SCALbx16_ARA0[9'd299] <= 33'h1ffffffff&-32'd4;
                   A_SINT_CC_SCALbx16_ARA0[9'd298] <= 33'h1ffffffff&32'd2;
                   A_SINT_CC_SCALbx16_ARA0[9'd297] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[9'd296] <= 33'h1ffffffff&-32'd1;
                   A_SINT_CC_SCALbx16_ARA0[9'd295] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[9'd294] <= 33'h1ffffffff&32'd6;
                   A_SINT_CC_SCALbx16_ARA0[9'd293] <= 33'h1ffffffff&32'd1;
                   A_SINT_CC_SCALbx16_ARA0[9'd292] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[9'd291] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[9'd290] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[9'd289] <= 33'h1ffffffff&-32'd3;
                   A_SINT_CC_SCALbx16_ARA0[9'd288] <= 33'h1ffffffff&32'd3;
                   A_SINT_CC_SCALbx16_ARA0[9'd287] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[9'd286] <= 33'h1ffffffff&32'd2;
                   A_SINT_CC_SCALbx16_ARA0[9'd285] <= 33'h1ffffffff&-32'd3;
                   A_SINT_CC_SCALbx16_ARA0[9'd284] <= 33'h1ffffffff&-32'd4;
                   A_SINT_CC_SCALbx16_ARA0[9'd283] <= 33'h1ffffffff&-32'd1;
                   A_SINT_CC_SCALbx16_ARA0[9'd282] <= 33'h1ffffffff&-32'd1;
                   A_SINT_CC_SCALbx16_ARA0[9'd281] <= 33'h1ffffffff&-32'd4;
                   A_SINT_CC_SCALbx16_ARA0[9'd280] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[9'd279] <= 33'h1ffffffff&-32'd4;
                   A_SINT_CC_SCALbx16_ARA0[9'd278] <= 33'h1ffffffff&-32'd5;
                   A_SINT_CC_SCALbx16_ARA0[9'd277] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[9'd276] <= 33'h1ffffffff&-32'd1;
                   A_SINT_CC_SCALbx16_ARA0[9'd275] <= 33'h1ffffffff&-32'd1;
                   A_SINT_CC_SCALbx16_ARA0[9'd274] <= 33'h1ffffffff&32'd1;
                   A_SINT_CC_SCALbx16_ARA0[9'd273] <= 33'h1ffffffff&32'd4;
                   A_SINT_CC_SCALbx16_ARA0[9'd272] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[9'd271] <= 33'h1ffffffff&32'd1;
                   A_SINT_CC_SCALbx16_ARA0[9'd270] <= 33'h1ffffffff&-32'd1;
                   A_SINT_CC_SCALbx16_ARA0[9'd269] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[9'd268] <= 33'h1ffffffff&32'd1;
                   A_SINT_CC_SCALbx16_ARA0[9'd267] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[9'd266] <= 33'h1ffffffff&32'd3;
                   A_SINT_CC_SCALbx16_ARA0[9'd265] <= 33'h1ffffffff&-32'd1;
                   A_SINT_CC_SCALbx16_ARA0[9'd264] <= 33'h1ffffffff&-32'd5;
                   A_SINT_CC_SCALbx16_ARA0[9'd263] <= 33'h1ffffffff&32'd2;
                   A_SINT_CC_SCALbx16_ARA0[9'd262] <= 33'h1ffffffff&32'd2;
                   A_SINT_CC_SCALbx16_ARA0[9'd261] <= 33'h1ffffffff&-32'd5;
                   A_SINT_CC_SCALbx16_ARA0[9'd260] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[9'd259] <= 33'h1ffffffff&-32'd5;
                   A_SINT_CC_SCALbx16_ARA0[9'd258] <= 33'h1ffffffff&-32'd6;
                   A_SINT_CC_SCALbx16_ARA0[9'd257] <= 33'h1ffffffff&-32'd1;
                   A_SINT_CC_SCALbx16_ARA0[9'd256] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[8'd255] <= 33'h1ffffffff&32'd1;
                   A_SINT_CC_SCALbx16_ARA0[8'd254] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[8'd253] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[8'd252] <= 33'h1ffffffff&32'd6;
                   A_SINT_CC_SCALbx16_ARA0[8'd251] <= 33'h1ffffffff&-32'd1;
                   A_SINT_CC_SCALbx16_ARA0[8'd250] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[8'd249] <= 33'h1ffffffff&-32'd3;
                   A_SINT_CC_SCALbx16_ARA0[8'd248] <= 33'h1ffffffff&-32'd1;
                   A_SINT_CC_SCALbx16_ARA0[8'd247] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[8'd246] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[8'd245] <= 33'h1ffffffff&-32'd1;
                   A_SINT_CC_SCALbx16_ARA0[8'd244] <= 33'h1ffffffff&-32'd5;
                   A_SINT_CC_SCALbx16_ARA0[8'd243] <= 33'h1ffffffff&-32'd1;
                   A_SINT_CC_SCALbx16_ARA0[8'd242] <= 33'h1ffffffff&-32'd1;
                   A_SINT_CC_SCALbx16_ARA0[8'd241] <= 33'h1ffffffff&-32'd3;
                   A_SINT_CC_SCALbx16_ARA0[8'd240] <= 33'h1ffffffff&32'd1;
                   A_SINT_CC_SCALbx16_ARA0[8'd239] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[8'd238] <= 33'h1ffffffff&-32'd4;
                   A_SINT_CC_SCALbx16_ARA0[8'd237] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[8'd236] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[8'd235] <= 33'h1ffffffff&32'd1;
                   A_SINT_CC_SCALbx16_ARA0[8'd234] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[8'd233] <= 33'h1ffffffff&32'd1;
                   A_SINT_CC_SCALbx16_ARA0[8'd232] <= 33'h1ffffffff&-32'd1;
                   A_SINT_CC_SCALbx16_ARA0[8'd231] <= 33'h1ffffffff&32'd2;
                   A_SINT_CC_SCALbx16_ARA0[8'd230] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[8'd229] <= 33'h1ffffffff&-32'd3;
                   A_SINT_CC_SCALbx16_ARA0[8'd228] <= 33'h1ffffffff&32'd1;
                   A_SINT_CC_SCALbx16_ARA0[8'd227] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[8'd226] <= 33'h1ffffffff&32'd2;
                   A_SINT_CC_SCALbx16_ARA0[8'd225] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[8'd224] <= 33'h1ffffffff&-32'd4;
                   A_SINT_CC_SCALbx16_ARA0[8'd223] <= 33'h1ffffffff&32'd1;
                   A_SINT_CC_SCALbx16_ARA0[8'd222] <= 33'h1ffffffff&32'd2;
                   A_SINT_CC_SCALbx16_ARA0[8'd221] <= 33'h1ffffffff&-32'd4;
                   A_SINT_CC_SCALbx16_ARA0[8'd220] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[8'd219] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[8'd218] <= 33'h1ffffffff&-32'd4;
                   A_SINT_CC_SCALbx16_ARA0[8'd217] <= 33'h1ffffffff&32'd2;
                   A_SINT_CC_SCALbx16_ARA0[8'd216] <= 33'h1ffffffff&-32'd1;
                   A_SINT_CC_SCALbx16_ARA0[8'd215] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[8'd214] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[8'd213] <= 33'h1ffffffff&-32'd1;
                   A_SINT_CC_SCALbx16_ARA0[8'd212] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[8'd211] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[8'd210] <= 33'h1ffffffff&32'd6;
                   A_SINT_CC_SCALbx16_ARA0[8'd209] <= 33'h1ffffffff&32'd4;
                   A_SINT_CC_SCALbx16_ARA0[8'd208] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[8'd207] <= 33'h1ffffffff&32'd2;
                   A_SINT_CC_SCALbx16_ARA0[8'd206] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[8'd205] <= 33'h1ffffffff&-32'd3;
                   A_SINT_CC_SCALbx16_ARA0[8'd204] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[8'd203] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[8'd202] <= 33'h1ffffffff&-32'd3;
                   A_SINT_CC_SCALbx16_ARA0[8'd201] <= 33'h1ffffffff&-32'd5;
                   A_SINT_CC_SCALbx16_ARA0[8'd200] <= 33'h1ffffffff&-32'd1;
                   A_SINT_CC_SCALbx16_ARA0[8'd199] <= 33'h1ffffffff&-32'd1;
                   A_SINT_CC_SCALbx16_ARA0[8'd198] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[8'd197] <= 33'h1ffffffff&32'd2;
                   A_SINT_CC_SCALbx16_ARA0[8'd196] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[8'd195] <= 33'h1ffffffff&-32'd3;
                   A_SINT_CC_SCALbx16_ARA0[8'd194] <= 33'h1ffffffff&-32'd3;
                   A_SINT_CC_SCALbx16_ARA0[8'd193] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[8'd192] <= 33'h1ffffffff&-32'd3;
                   A_SINT_CC_SCALbx16_ARA0[8'd191] <= 33'h1ffffffff&-32'd3;
                   A_SINT_CC_SCALbx16_ARA0[8'd190] <= 33'h1ffffffff&32'd4;
                   A_SINT_CC_SCALbx16_ARA0[8'd189] <= 33'h1ffffffff&32'd6;
                   A_SINT_CC_SCALbx16_ARA0[8'd188] <= 33'h1ffffffff&-32'd3;
                   A_SINT_CC_SCALbx16_ARA0[8'd187] <= 33'h1ffffffff&32'd2;
                   A_SINT_CC_SCALbx16_ARA0[8'd186] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[8'd185] <= 33'h1ffffffff&-32'd4;
                   A_SINT_CC_SCALbx16_ARA0[8'd184] <= 33'h1ffffffff&32'd2;
                   A_SINT_CC_SCALbx16_ARA0[8'd183] <= 33'h1ffffffff&-32'd3;
                   A_SINT_CC_SCALbx16_ARA0[8'd182] <= 33'h1ffffffff&-32'd4;
                   A_SINT_CC_SCALbx16_ARA0[8'd181] <= 33'h1ffffffff&-32'd6;
                   A_SINT_CC_SCALbx16_ARA0[8'd180] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[8'd179] <= 33'h1ffffffff&-32'd4;
                   A_SINT_CC_SCALbx16_ARA0[8'd178] <= 33'h1ffffffff&-32'd3;
                   A_SINT_CC_SCALbx16_ARA0[8'd177] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[8'd176] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[8'd175] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[8'd174] <= 33'h1ffffffff&32'd3;
                   A_SINT_CC_SCALbx16_ARA0[8'd173] <= 33'h1ffffffff&32'd1;
                   A_SINT_CC_SCALbx16_ARA0[8'd172] <= 33'h1ffffffff&-32'd1;
                   A_SINT_CC_SCALbx16_ARA0[8'd171] <= 33'h1ffffffff&32'd1;
                   A_SINT_CC_SCALbx16_ARA0[8'd170] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[8'd169] <= 33'h1ffffffff&-32'd3;
                   A_SINT_CC_SCALbx16_ARA0[8'd168] <= 33'h1ffffffff&32'd5;
                   A_SINT_CC_SCALbx16_ARA0[8'd167] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[8'd166] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[8'd165] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[8'd164] <= 33'h1ffffffff&-32'd5;
                   A_SINT_CC_SCALbx16_ARA0[8'd163] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[8'd162] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[8'd161] <= 33'h1ffffffff&-32'd5;
                   A_SINT_CC_SCALbx16_ARA0[8'd160] <= 33'h1ffffffff&-32'd1;
                   A_SINT_CC_SCALbx16_ARA0[8'd159] <= 33'h1ffffffff&-32'd1;
                   A_SINT_CC_SCALbx16_ARA0[8'd158] <= 33'h1ffffffff&-32'd5;
                   A_SINT_CC_SCALbx16_ARA0[8'd157] <= 33'h1ffffffff&32'd4;
                   A_SINT_CC_SCALbx16_ARA0[8'd156] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[8'd155] <= 33'h1ffffffff&-32'd1;
                   A_SINT_CC_SCALbx16_ARA0[8'd154] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[8'd153] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[8'd152] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[8'd151] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[8'd150] <= 33'h1ffffffff&32'd2;
                   A_SINT_CC_SCALbx16_ARA0[8'd149] <= 33'h1ffffffff&32'd2;
                   A_SINT_CC_SCALbx16_ARA0[8'd148] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[8'd147] <= 33'h1ffffffff&32'd5;
                   A_SINT_CC_SCALbx16_ARA0[8'd146] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[8'd145] <= 33'h1ffffffff&-32'd3;
                   A_SINT_CC_SCALbx16_ARA0[8'd144] <= 33'h1ffffffff&32'd1;
                   A_SINT_CC_SCALbx16_ARA0[8'd143] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[8'd142] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[8'd141] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[8'd140] <= 33'h1ffffffff&-32'd1;
                   A_SINT_CC_SCALbx16_ARA0[8'd139] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[8'd138] <= 33'h1ffffffff&-32'd3;
                   A_SINT_CC_SCALbx16_ARA0[8'd137] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[8'd136] <= 33'h1ffffffff&-32'd1;
                   A_SINT_CC_SCALbx16_ARA0[8'd135] <= 33'h1ffffffff&-32'd1;
                   A_SINT_CC_SCALbx16_ARA0[8'd134] <= 33'h1ffffffff&32'd2;
                   A_SINT_CC_SCALbx16_ARA0[8'd133] <= 33'h1ffffffff&32'd3;
                   A_SINT_CC_SCALbx16_ARA0[8'd132] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[8'd131] <= 33'h1ffffffff&32'd2;
                   A_SINT_CC_SCALbx16_ARA0[8'd130] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[8'd129] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[8'd128] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[7'd127] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[7'd126] <= 33'h1ffffffff&32'd6;
                   A_SINT_CC_SCALbx16_ARA0[7'd125] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[7'd124] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[7'd123] <= 33'h1ffffffff&32'd1;
                   A_SINT_CC_SCALbx16_ARA0[7'd122] <= 33'h1ffffffff&32'd1;
                   A_SINT_CC_SCALbx16_ARA0[7'd121] <= 33'h1ffffffff&-32'd3;
                   A_SINT_CC_SCALbx16_ARA0[7'd120] <= 33'h1ffffffff&-32'd1;
                   A_SINT_CC_SCALbx16_ARA0[7'd119] <= 33'h1ffffffff&-32'd5;
                   A_SINT_CC_SCALbx16_ARA0[7'd118] <= 33'h1ffffffff&-32'd7;
                   A_SINT_CC_SCALbx16_ARA0[7'd117] <= 33'h1ffffffff&-32'd1;
                   A_SINT_CC_SCALbx16_ARA0[7'd116] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[7'd115] <= 33'h1ffffffff&32'd1;
                   A_SINT_CC_SCALbx16_ARA0[7'd114] <= 33'h1ffffffff&-32'd3;
                   A_SINT_CC_SCALbx16_ARA0[7'd113] <= 33'h1ffffffff&-32'd1;
                   A_SINT_CC_SCALbx16_ARA0[7'd112] <= 33'h1ffffffff&-32'd1;
                   A_SINT_CC_SCALbx16_ARA0[7'd111] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[7'd110] <= 33'h1ffffffff&-32'd3;
                   A_SINT_CC_SCALbx16_ARA0[7'd109] <= 33'h1ffffffff&-32'd4;
                   A_SINT_CC_SCALbx16_ARA0[7'd108] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[7'd107] <= 33'h1ffffffff&-32'd3;
                   A_SINT_CC_SCALbx16_ARA0[7'd106] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[7'd105] <= 33'h1ffffffff&32'd5;
                   A_SINT_CC_SCALbx16_ARA0[7'd104] <= 33'h1ffffffff&-32'd5;
                   A_SINT_CC_SCALbx16_ARA0[7'd103] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[7'd102] <= 33'h1ffffffff&32'd1;
                   A_SINT_CC_SCALbx16_ARA0[7'd101] <= 33'h1ffffffff&-32'd3;
                   A_SINT_CC_SCALbx16_ARA0[7'd100] <= 33'h1ffffffff&32'd1;
                   A_SINT_CC_SCALbx16_ARA0[7'd99] <= 33'h1ffffffff&32'd7;
                   A_SINT_CC_SCALbx16_ARA0[7'd98] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[7'd97] <= 33'h1ffffffff&-32'd1;
                   A_SINT_CC_SCALbx16_ARA0[7'd96] <= 33'h1ffffffff&-32'd3;
                   A_SINT_CC_SCALbx16_ARA0[7'd95] <= 33'h1ffffffff&-32'd3;
                   A_SINT_CC_SCALbx16_ARA0[7'd94] <= 33'h1ffffffff&-32'd4;
                   A_SINT_CC_SCALbx16_ARA0[7'd93] <= 33'h1ffffffff&-32'd5;
                   A_SINT_CC_SCALbx16_ARA0[7'd92] <= 33'h1ffffffff&-32'd5;
                   A_SINT_CC_SCALbx16_ARA0[7'd91] <= 33'h1ffffffff&-32'd4;
                   A_SINT_CC_SCALbx16_ARA0[7'd90] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[7'd89] <= 33'h1ffffffff&32'd2;
                   A_SINT_CC_SCALbx16_ARA0[7'd88] <= 33'h1ffffffff&-32'd5;
                   A_SINT_CC_SCALbx16_ARA0[7'd87] <= 33'h1ffffffff&32'd1;
                   A_SINT_CC_SCALbx16_ARA0[7'd86] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[7'd85] <= 33'h1ffffffff&-32'd5;
                   A_SINT_CC_SCALbx16_ARA0[7'd84] <= 33'h1ffffffff&32'd9;
                   A_SINT_CC_SCALbx16_ARA0[7'd83] <= 33'h1ffffffff&-32'd5;
                   A_SINT_CC_SCALbx16_ARA0[7'd82] <= 33'h1ffffffff&-32'd6;
                   A_SINT_CC_SCALbx16_ARA0[7'd81] <= 33'h1ffffffff&-32'd4;
                   A_SINT_CC_SCALbx16_ARA0[7'd80] <= 33'h1ffffffff&-32'd4;
                   A_SINT_CC_SCALbx16_ARA0[7'd79] <= 33'h1ffffffff&-32'd4;
                   A_SINT_CC_SCALbx16_ARA0[7'd78] <= 33'h1ffffffff&-32'd7;
                   A_SINT_CC_SCALbx16_ARA0[7'd77] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[7'd76] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[7'd75] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[7'd74] <= 33'h1ffffffff&-32'd1;
                   A_SINT_CC_SCALbx16_ARA0[7'd73] <= 33'h1ffffffff&32'd2;
                   A_SINT_CC_SCALbx16_ARA0[7'd72] <= 33'h1ffffffff&-32'd1;
                   A_SINT_CC_SCALbx16_ARA0[7'd71] <= 33'h1ffffffff&32'd1;
                   A_SINT_CC_SCALbx16_ARA0[7'd70] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[7'd69] <= 33'h1ffffffff&-32'd3;
                   A_SINT_CC_SCALbx16_ARA0[7'd68] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[7'd67] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[7'd66] <= 33'h1ffffffff&32'd1;
                   A_SINT_CC_SCALbx16_ARA0[7'd65] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[7'd64] <= 33'h1ffffffff&-32'd5;
                   A_SINT_CC_SCALbx16_ARA0[6'd63] <= 33'h1ffffffff&32'd4;
                   A_SINT_CC_SCALbx16_ARA0[6'd62] <= 33'h1ffffffff&32'd3;
                   A_SINT_CC_SCALbx16_ARA0[6'd61] <= 33'h1ffffffff&-32'd5;
                   A_SINT_CC_SCALbx16_ARA0[6'd60] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[6'd59] <= 33'h1ffffffff&-32'd4;
                   A_SINT_CC_SCALbx16_ARA0[6'd58] <= 33'h1ffffffff&-32'd7;
                   A_SINT_CC_SCALbx16_ARA0[6'd57] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[6'd56] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[6'd55] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[6'd54] <= 33'h1ffffffff&-32'd1;
                   A_SINT_CC_SCALbx16_ARA0[6'd53] <= 33'h1ffffffff&32'd2;
                   A_SINT_CC_SCALbx16_ARA0[6'd52] <= 33'h1ffffffff&-32'd1;
                   A_SINT_CC_SCALbx16_ARA0[6'd51] <= 33'h1ffffffff&32'd2;
                   A_SINT_CC_SCALbx16_ARA0[6'd50] <= 33'h1ffffffff&-32'd3;
                   A_SINT_CC_SCALbx16_ARA0[6'd49] <= 33'h1ffffffff&-32'd4;
                   A_SINT_CC_SCALbx16_ARA0[6'd48] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[6'd47] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[6'd46] <= 33'h1ffffffff&32'd1;
                   A_SINT_CC_SCALbx16_ARA0[6'd45] <= 33'h1ffffffff&32'd1;
                   A_SINT_CC_SCALbx16_ARA0[6'd44] <= 33'h1ffffffff&-32'd6;
                   A_SINT_CC_SCALbx16_ARA0[6'd43] <= 33'h1ffffffff&32'd3;
                   A_SINT_CC_SCALbx16_ARA0[6'd42] <= 33'h1ffffffff&32'd4;
                   A_SINT_CC_SCALbx16_ARA0[6'd41] <= 33'h1ffffffff&-32'd5;
                   A_SINT_CC_SCALbx16_ARA0[6'd40] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[6'd39] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[6'd38] <= 33'h1ffffffff&-32'd8;
                   A_SINT_CC_SCALbx16_ARA0[6'd37] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[6'd36] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[6'd35] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[6'd34] <= 33'h1ffffffff&-32'd4;
                   A_SINT_CC_SCALbx16_ARA0[6'd33] <= 33'h1ffffffff&-32'd5;
                   A_SINT_CC_SCALbx16_ARA0[6'd32] <= 33'h1ffffffff&-32'd3;
                   A_SINT_CC_SCALbx16_ARA0[5'd31] <= 33'h1ffffffff&-32'd4;
                   A_SINT_CC_SCALbx16_ARA0[5'd30] <= 33'h1ffffffff&-32'd5;
                   A_SINT_CC_SCALbx16_ARA0[5'd29] <= 33'h1ffffffff&-32'd6;
                   A_SINT_CC_SCALbx16_ARA0[5'd28] <= 33'h1ffffffff&-32'd5;
                   A_SINT_CC_SCALbx16_ARA0[5'd27] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[5'd26] <= 33'h1ffffffff&-32'd3;
                   A_SINT_CC_SCALbx16_ARA0[5'd25] <= 33'h1ffffffff&-32'd3;
                   A_SINT_CC_SCALbx16_ARA0[5'd24] <= 33'h1ffffffff&-32'd4;
                   A_SINT_CC_SCALbx16_ARA0[5'd23] <= 33'h1ffffffff&-32'd5;
                   A_SINT_CC_SCALbx16_ARA0[5'd22] <= 33'h1ffffffff&-32'd5;
                   A_SINT_CC_SCALbx16_ARA0[5'd21] <= 33'h1ffffffff&32'd12;
                   A_SINT_CC_SCALbx16_ARA0[5'd20] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[5'd19] <= 33'h1ffffffff&-32'd3;
                   A_SINT_CC_SCALbx16_ARA0[5'd18] <= 33'h1ffffffff&-32'd1;
                   A_SINT_CC_SCALbx16_ARA0[5'd17] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[5'd16] <= 33'h1ffffffff&32'd1;
                   A_SINT_CC_SCALbx16_ARA0[4'd15] <= 33'h1ffffffff&32'd1;
                   A_SINT_CC_SCALbx16_ARA0[4'd14] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[4'd13] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[4'd12] <= 33'h1ffffffff&32'd1;
                   A_SINT_CC_SCALbx16_ARA0[4'd11] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[4'd10] <= 33'h1ffffffff&-32'd1;
                   A_SINT_CC_SCALbx16_ARA0[4'd9] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[4'd8] <= 33'h1ffffffff&-32'd1;
                   A_SINT_CC_SCALbx16_ARA0[3'd7] <= 33'h1ffffffff&-32'd1;
                   A_SINT_CC_SCALbx16_ARA0[3'd6] <= 33'h1ffffffff&-32'd1;
                   A_SINT_CC_SCALbx16_ARA0[3'd5] <= 33'h1ffffffff&32'd1;
                   A_SINT_CC_SCALbx16_ARA0[3'd4] <= 33'h1ffffffff&-32'd4;
                   A_SINT_CC_SCALbx16_ARA0[2'd3] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[2'd2] <= 33'h1ffffffff&32'd0;
                   A_SINT_CC_SCALbx16_ARA0[1'd1] <= 33'h1ffffffff&-32'd2;
                   A_SINT_CC_SCALbx16_ARA0[0] <= 33'h1ffffffff&32'd2;
                   A_16_SS_CC_SCALbx10_ARA0[7'd74] <= 17'h1ffff&16'd108;
                   A_16_SS_CC_SCALbx10_ARA0[7'd73] <= 17'h1ffff&16'd112;
                   A_16_SS_CC_SCALbx10_ARA0[7'd72] <= 17'h1ffff&16'd105;
                   A_16_SS_CC_SCALbx10_ARA0[7'd71] <= 17'h1ffff&16'd116;
                   A_16_SS_CC_SCALbx10_ARA0[7'd70] <= 17'h1ffff&16'd101;
                   A_16_SS_CC_SCALbx10_ARA0[7'd69] <= 17'h1ffff&16'd121;
                   A_16_SS_CC_SCALbx10_ARA0[7'd68] <= 17'h1ffff&16'd103;
                   A_16_SS_CC_SCALbx10_ARA0[7'd67] <= 17'h1ffff&16'd113;
                   A_16_SS_CC_SCALbx10_ARA0[7'd66] <= 17'h1ffff&16'd105;
                   A_16_SS_CC_SCALbx10_ARA0[7'd65] <= 17'h1ffff&16'd114;
                   A_16_SS_CC_SCALbx10_ARA0[7'd64] <= 17'h1ffff&16'd97;
                   A_16_SS_CC_SCALbx10_ARA0[6'd63] <= 17'h1ffff&16'd118;
                   A_16_SS_CC_SCALbx10_ARA0[6'd62] <= 17'h1ffff&16'd101;
                   A_16_SS_CC_SCALbx10_ARA0[6'd61] <= 17'h1ffff&16'd101;
                   A_16_SS_CC_SCALbx10_ARA0[6'd60] <= 17'h1ffff&16'd118;
                   A_16_SS_CC_SCALbx10_ARA0[6'd59] <= 17'h1ffff&16'd108;
                   A_16_SS_CC_SCALbx10_ARA0[6'd58] <= 17'h1ffff&16'd100;
                   A_16_SS_CC_SCALbx10_ARA0[6'd57] <= 17'h1ffff&16'd101;
                   A_16_SS_CC_SCALbx10_ARA0[6'd56] <= 17'h1ffff&16'd101;
                   A_16_SS_CC_SCALbx10_ARA0[6'd55] <= 17'h1ffff&16'd108;
                   A_16_SS_CC_SCALbx10_ARA0[6'd54] <= 17'h1ffff&16'd114;
                   A_16_SS_CC_SCALbx10_ARA0[6'd53] <= 17'h1ffff&16'd108;
                   A_16_SS_CC_SCALbx10_ARA0[6'd52] <= 17'h1ffff&16'd100;
                   A_16_SS_CC_SCALbx10_ARA0[6'd51] <= 17'h1ffff&16'd108;
                   A_16_SS_CC_SCALbx10_ARA0[6'd50] <= 17'h1ffff&16'd114;
                   A_16_SS_CC_SCALbx10_ARA0[6'd49] <= 17'h1ffff&16'd104;
                   A_16_SS_CC_SCALbx10_ARA0[6'd48] <= 17'h1ffff&16'd115;
                   A_16_SS_CC_SCALbx10_ARA0[6'd47] <= 17'h1ffff&16'd112;
                   A_16_SS_CC_SCALbx10_ARA0[6'd46] <= 17'h1ffff&16'd112;
                   A_16_SS_CC_SCALbx10_ARA0[6'd45] <= 17'h1ffff&16'd116;
                   A_16_SS_CC_SCALbx10_ARA0[6'd44] <= 17'h1ffff&16'd118;
                   A_16_SS_CC_SCALbx10_ARA0[6'd43] <= 17'h1ffff&16'd114;
                   A_16_SS_CC_SCALbx10_ARA0[6'd42] <= 17'h1ffff&16'd121;
                   A_16_SS_CC_SCALbx10_ARA0[6'd41] <= 17'h1ffff&16'd116;
                   A_16_SS_CC_SCALbx10_ARA0[6'd40] <= 17'h1ffff&16'd112;
                   A_16_SS_CC_SCALbx10_ARA0[6'd39] <= 17'h1ffff&16'd103;
                   A_16_SS_CC_SCALbx10_ARA0[6'd38] <= 17'h1ffff&16'd101;
                   A_16_SS_CC_SCALbx10_ARA0[6'd37] <= 17'h1ffff&16'd103;
                   A_16_SS_CC_SCALbx10_ARA0[6'd36] <= 17'h1ffff&16'd101;
                   A_16_SS_CC_SCALbx10_ARA0[6'd35] <= 17'h1ffff&16'd118;
                   A_16_SS_CC_SCALbx10_ARA0[6'd34] <= 17'h1ffff&16'd114;
                   A_16_SS_CC_SCALbx10_ARA0[6'd33] <= 17'h1ffff&16'd99;
                   A_16_SS_CC_SCALbx10_ARA0[6'd32] <= 17'h1ffff&16'd103;
                   A_16_SS_CC_SCALbx10_ARA0[5'd31] <= 17'h1ffff&16'd108;
                   A_16_SS_CC_SCALbx10_ARA0[5'd30] <= 17'h1ffff&16'd114;
                   A_16_SS_CC_SCALbx10_ARA0[5'd29] <= 17'h1ffff&16'd107;
                   A_16_SS_CC_SCALbx10_ARA0[5'd28] <= 17'h1ffff&16'd108;
                   A_16_SS_CC_SCALbx10_ARA0[5'd27] <= 17'h1ffff&16'd105;
                   A_16_SS_CC_SCALbx10_ARA0[5'd26] <= 17'h1ffff&16'd97;
                   A_16_SS_CC_SCALbx10_ARA0[5'd25] <= 17'h1ffff&16'd105;
                   A_16_SS_CC_SCALbx10_ARA0[5'd24] <= 17'h1ffff&16'd113;
                   A_16_SS_CC_SCALbx10_ARA0[5'd23] <= 17'h1ffff&16'd101;
                   A_16_SS_CC_SCALbx10_ARA0[5'd22] <= 17'h1ffff&16'd97;
                   A_16_SS_CC_SCALbx10_ARA0[5'd21] <= 17'h1ffff&16'd101;
                   A_16_SS_CC_SCALbx10_ARA0[5'd20] <= 17'h1ffff&16'd112;
                   A_16_SS_CC_SCALbx10_ARA0[5'd19] <= 17'h1ffff&16'd121;
                   A_16_SS_CC_SCALbx10_ARA0[5'd18] <= 17'h1ffff&16'd115;
                   A_16_SS_CC_SCALbx10_ARA0[5'd17] <= 17'h1ffff&16'd116;
                   A_16_SS_CC_SCALbx10_ARA0[5'd16] <= 17'h1ffff&16'd103;
                   A_16_SS_CC_SCALbx10_ARA0[4'd15] <= 17'h1ffff&16'd108;
                   A_16_SS_CC_SCALbx10_ARA0[4'd14] <= 17'h1ffff&16'd108;
                   A_16_SS_CC_SCALbx10_ARA0[4'd13] <= 17'h1ffff&16'd114;
                   A_16_SS_CC_SCALbx10_ARA0[4'd12] <= 17'h1ffff&16'd110;
                   A_16_SS_CC_SCALbx10_ARA0[4'd11] <= 17'h1ffff&16'd97;
                   A_16_SS_CC_SCALbx10_ARA0[4'd10] <= 17'h1ffff&16'd121;
                   A_16_SS_CC_SCALbx10_ARA0[4'd9] <= 17'h1ffff&16'd101;
                   A_16_SS_CC_SCALbx10_ARA0[4'd8] <= 17'h1ffff&16'd112;
                   A_16_SS_CC_SCALbx10_ARA0[3'd7] <= 17'h1ffff&16'd114;
                   A_16_SS_CC_SCALbx10_ARA0[3'd6] <= 17'h1ffff&16'd102;
                   A_16_SS_CC_SCALbx10_ARA0[3'd5] <= 17'h1ffff&16'd112;
                   A_16_SS_CC_SCALbx10_ARA0[3'd4] <= 17'h1ffff&16'd105;
                   A_16_SS_CC_SCALbx10_ARA0[2'd3] <= 17'h1ffff&16'd97;
                   A_16_SS_CC_SCALbx10_ARA0[2'd2] <= 17'h1ffff&16'd101;
                   A_16_SS_CC_SCALbx10_ARA0[1'd1] <= 17'h1ffff&16'd112;
                   A_16_SS_CC_SCALbx10_ARA0[0] <= 17'h1ffff&16'd112;
                   A_16_SS_CC_SCALbx14_ARC0[7'd76] <= 17'h1ffff&16'd110;
                   A_16_SS_CC_SCALbx14_ARC0[7'd75] <= 17'h1ffff&16'd101;
                   A_16_SS_CC_SCALbx14_ARC0[7'd74] <= 17'h1ffff&16'd113;
                   A_16_SS_CC_SCALbx14_ARC0[7'd73] <= 17'h1ffff&16'd114;
                   A_16_SS_CC_SCALbx14_ARC0[7'd72] <= 17'h1ffff&16'd118;
                   A_16_SS_CC_SCALbx14_ARC0[7'd71] <= 17'h1ffff&16'd101;
                   A_16_SS_CC_SCALbx14_ARC0[7'd70] <= 17'h1ffff&16'd107;
                   A_16_SS_CC_SCALbx14_ARC0[7'd69] <= 17'h1ffff&16'd97;
                   A_16_SS_CC_SCALbx14_ARC0[7'd68] <= 17'h1ffff&16'd101;
                   A_16_SS_CC_SCALbx14_ARC0[7'd67] <= 17'h1ffff&16'd101;
                   A_16_SS_CC_SCALbx14_ARC0[7'd66] <= 17'h1ffff&16'd108;
                   A_16_SS_CC_SCALbx14_ARC0[7'd65] <= 17'h1ffff&16'd97;
                   A_16_SS_CC_SCALbx14_ARC0[7'd64] <= 17'h1ffff&16'd101;
                   A_16_SS_CC_SCALbx14_ARC0[6'd63] <= 17'h1ffff&16'd113;
                   A_16_SS_CC_SCALbx14_ARC0[6'd62] <= 17'h1ffff&16'd115;
                   A_16_SS_CC_SCALbx14_ARC0[6'd61] <= 17'h1ffff&16'd103;
                   A_16_SS_CC_SCALbx14_ARC0[6'd60] <= 17'h1ffff&16'd119;
                   A_16_SS_CC_SCALbx14_ARC0[6'd59] <= 17'h1ffff&16'd118;
                   A_16_SS_CC_SCALbx14_ARC0[6'd58] <= 17'h1ffff&16'd101;
                   A_16_SS_CC_SCALbx14_ARC0[6'd57] <= 17'h1ffff&16'd108;
                   A_16_SS_CC_SCALbx14_ARC0[6'd56] <= 17'h1ffff&16'd115;
                   A_16_SS_CC_SCALbx14_ARC0[6'd55] <= 17'h1ffff&16'd114;
                   A_16_SS_CC_SCALbx14_ARC0[6'd54] <= 17'h1ffff&16'd107;
                   A_16_SS_CC_SCALbx14_ARC0[6'd53] <= 17'h1ffff&16'd118;
                   A_16_SS_CC_SCALbx14_ARC0[6'd52] <= 17'h1ffff&16'd105;
                   A_16_SS_CC_SCALbx14_ARC0[6'd51] <= 17'h1ffff&16'd113;
                   A_16_SS_CC_SCALbx14_ARC0[6'd50] <= 17'h1ffff&16'd108;
                   A_16_SS_CC_SCALbx14_ARC0[6'd49] <= 17'h1ffff&16'd107;
                   A_16_SS_CC_SCALbx14_ARC0[6'd48] <= 17'h1ffff&16'd108;
                   A_16_SS_CC_SCALbx14_ARC0[6'd47] <= 17'h1ffff&16'd121;
                   A_16_SS_CC_SCALbx14_ARC0[6'd46] <= 17'h1ffff&16'd108;
                   A_16_SS_CC_SCALbx14_ARC0[6'd45] <= 17'h1ffff&16'd107;
                   A_16_SS_CC_SCALbx14_ARC0[6'd44] <= 17'h1ffff&16'd109;
                   A_16_SS_CC_SCALbx14_ARC0[6'd43] <= 17'h1ffff&16'd100;
                   A_16_SS_CC_SCALbx14_ARC0[6'd42] <= 17'h1ffff&16'd103;
                   A_16_SS_CC_SCALbx14_ARC0[6'd41] <= 17'h1ffff&16'd119;
                   A_16_SS_CC_SCALbx14_ARC0[6'd40] <= 17'h1ffff&16'd113;
                   A_16_SS_CC_SCALbx14_ARC0[6'd39] <= 17'h1ffff&16'd115;
                   A_16_SS_CC_SCALbx14_ARC0[6'd38] <= 17'h1ffff&16'd104;
                   A_16_SS_CC_SCALbx14_ARC0[6'd37] <= 17'h1ffff&16'd104;
                   A_16_SS_CC_SCALbx14_ARC0[6'd36] <= 17'h1ffff&16'd112;
                   A_16_SS_CC_SCALbx14_ARC0[6'd35] <= 17'h1ffff&16'd110;
                   A_16_SS_CC_SCALbx14_ARC0[6'd34] <= 17'h1ffff&16'd107;
                   A_16_SS_CC_SCALbx14_ARC0[6'd33] <= 17'h1ffff&16'd107;
                   A_16_SS_CC_SCALbx14_ARC0[6'd32] <= 17'h1ffff&16'd118;
                   A_16_SS_CC_SCALbx14_ARC0[5'd31] <= 17'h1ffff&16'd105;
                   A_16_SS_CC_SCALbx14_ARC0[5'd30] <= 17'h1ffff&16'd102;
                   A_16_SS_CC_SCALbx14_ARC0[5'd29] <= 17'h1ffff&16'd107;
                   A_16_SS_CC_SCALbx14_ARC0[5'd28] <= 17'h1ffff&16'd108;
                   A_16_SS_CC_SCALbx14_ARC0[5'd27] <= 17'h1ffff&16'd112;
                   A_16_SS_CC_SCALbx14_ARC0[5'd26] <= 17'h1ffff&16'd112;
                   A_16_SS_CC_SCALbx14_ARC0[5'd25] <= 17'h1ffff&16'd101;
                   A_16_SS_CC_SCALbx14_ARC0[5'd24] <= 17'h1ffff&16'd114;
                   A_16_SS_CC_SCALbx14_ARC0[5'd23] <= 17'h1ffff&16'd107;
                   A_16_SS_CC_SCALbx14_ARC0[5'd22] <= 17'h1ffff&16'd101;
                   A_16_SS_CC_SCALbx14_ARC0[5'd21] <= 17'h1ffff&16'd108;
                   A_16_SS_CC_SCALbx14_ARC0[5'd20] <= 17'h1ffff&16'd100;
                   A_16_SS_CC_SCALbx14_ARC0[5'd19] <= 17'h1ffff&16'd99;
                   A_16_SS_CC_SCALbx14_ARC0[5'd18] <= 17'h1ffff&16'd100;
                   A_16_SS_CC_SCALbx14_ARC0[5'd17] <= 17'h1ffff&16'd107;
                   A_16_SS_CC_SCALbx14_ARC0[5'd16] <= 17'h1ffff&16'd108;
                   A_16_SS_CC_SCALbx14_ARC0[4'd15] <= 17'h1ffff&16'd108;
                   A_16_SS_CC_SCALbx14_ARC0[4'd14] <= 17'h1ffff&16'd121;
                   A_16_SS_CC_SCALbx14_ARC0[4'd13] <= 17'h1ffff&16'd101;
                   A_16_SS_CC_SCALbx14_ARC0[4'd12] <= 17'h1ffff&16'd113;
                   A_16_SS_CC_SCALbx14_ARC0[4'd11] <= 17'h1ffff&16'd107;
                   A_16_SS_CC_SCALbx14_ARC0[4'd10] <= 17'h1ffff&16'd97;
                   A_16_SS_CC_SCALbx14_ARC0[4'd9] <= 17'h1ffff&16'd101;
                   A_16_SS_CC_SCALbx14_ARC0[4'd8] <= 17'h1ffff&16'd116;
                   A_16_SS_CC_SCALbx14_ARC0[3'd7] <= 17'h1ffff&16'd107;
                   A_16_SS_CC_SCALbx14_ARC0[3'd6] <= 17'h1ffff&16'd116;
                   A_16_SS_CC_SCALbx14_ARC0[3'd5] <= 17'h1ffff&16'd105;
                   A_16_SS_CC_SCALbx14_ARC0[3'd4] <= 17'h1ffff&16'd108;
                   A_16_SS_CC_SCALbx14_ARC0[2'd3] <= 17'h1ffff&16'd107;
                   A_16_SS_CC_SCALbx14_ARC0[2'd2] <= 17'h1ffff&16'd104;
                   A_16_SS_CC_SCALbx14_ARC0[1'd1] <= 17'h1ffff&16'd107;
                   A_16_SS_CC_SCALbx14_ARC0[0] <= 17'h1ffff&16'd100;
                   A_16_SS_CC_SCALbx12_ARB0[5'd19] <= 17'h1ffff&16'd121;
                   A_16_SS_CC_SCALbx12_ARB0[5'd18] <= 17'h1ffff&16'd119;
                   A_16_SS_CC_SCALbx12_ARB0[5'd17] <= 17'h1ffff&16'd118;
                   A_16_SS_CC_SCALbx12_ARB0[5'd16] <= 17'h1ffff&16'd116;
                   A_16_SS_CC_SCALbx12_ARB0[4'd15] <= 17'h1ffff&16'd115;
                   A_16_SS_CC_SCALbx12_ARB0[4'd14] <= 17'h1ffff&16'd114;
                   A_16_SS_CC_SCALbx12_ARB0[4'd13] <= 17'h1ffff&16'd113;
                   A_16_SS_CC_SCALbx12_ARB0[4'd12] <= 17'h1ffff&16'd112;
                   A_16_SS_CC_SCALbx12_ARB0[4'd11] <= 17'h1ffff&16'd110;
                   A_16_SS_CC_SCALbx12_ARB0[4'd10] <= 17'h1ffff&16'd109;
                   A_16_SS_CC_SCALbx12_ARB0[4'd9] <= 17'h1ffff&16'd108;
                   A_16_SS_CC_SCALbx12_ARB0[4'd8] <= 17'h1ffff&16'd107;
                   A_16_SS_CC_SCALbx12_ARB0[3'd7] <= 17'h1ffff&16'd105;
                   A_16_SS_CC_SCALbx12_ARB0[3'd6] <= 17'h1ffff&16'd104;
                   A_16_SS_CC_SCALbx12_ARB0[3'd5] <= 17'h1ffff&16'd103;
                   A_16_SS_CC_SCALbx12_ARB0[3'd4] <= 17'h1ffff&16'd102;
                   A_16_SS_CC_SCALbx12_ARB0[2'd3] <= 17'h1ffff&16'd101;
                   A_16_SS_CC_SCALbx12_ARB0[2'd2] <= 17'h1ffff&16'd100;
                   A_16_SS_CC_SCALbx12_ARB0[1'd1] <= 17'h1ffff&16'd99;
                   A_16_SS_CC_SCALbx12_ARB0[0] <= 17'h1ffff&16'd97;
                   end 
                  
              2'd3/*3:US*/: if (((33'h1ffffffff&32'd1+TSPin0_6_V_0)<(33'h1ffffffff&32'h4d)))  begin 
                       xpc10 <= 6'd41/*41:xpc10:41*/;
                       TSPen1_8_V_0 <= 33'h1ffffffff&32'd0;
                       TSPin0_6_V_0 <= 33'h1ffffffff&32'd1+TSPin0_6_V_0;
                       A_SINT_CC_SCALbx26_ARJ0[TSPin0_6_V_0] <= 33'h1ffffffff&TSPe1_SPILL_256;
                       end 
                       else  begin 
                       xpc10 <= 3'd4/*4:xpc10:4*/;
                       TSPru0_12_V_0 <= 33'h1ffffffff&32'd0;
                       phase <= 33'h1ffffffff&32'd3;
                       TSPin0_6_V_0 <= 33'h1ffffffff&32'd1+TSPin0_6_V_0;
                       A_SINT_CC_SCALbx26_ARJ0[TSPin0_6_V_0] <= 33'h1ffffffff&TSPe1_SPILL_256;
                       end 
                      
              3'd4/*4:US*/: if ((TSPru0_12_V_0<(33'h1ffffffff&32'd1)))  xpc10 <= 5'd16/*16:xpc10:16*/;
                   else  begin 
                       xpc10 <= 3'd5/*5:xpc10:5*/;
                       A_UINT_CC_SCALbx38_crc_reg <= 33'h1ffffffff&-32'd1;
                       phase <= 33'h1ffffffff&32'd12;
                       end 
                      
              5'd19/*19:US*/: if ((TSPru0_12_V_1<2'd3))  begin 
                       xpc10 <= 5'd20/*20:xpc10:20*/;
                       TSPen0_17_V_0 <= 33'h1ffffffff&32'd0;
                       TSPne2_10_V_1 <= 33'h1ffffffff&((32'd1+TSPru0_12_V_1)%2'd2);
                       TSPne2_10_V_0 <= 33'h1ffffffff&(TSPru0_12_V_1%2'd2);
                       phase <= 33'h1ffffffff&32'd4;
                       end 
                       else  begin 
                       xpc10 <= 3'd4/*4:xpc10:4*/;
                       TSPru0_12_V_0 <= 33'h1ffffffff&32'd1+TSPru0_12_V_0;
                       end 
                      
              5'd22/*22:US*/: if ((TSPne2_10_V_3<(33'h1ffffffff&32'h4d)))  xpc10 <= 6'd32/*32:xpc10:32*/;
                   else  begin 
                       xpc10 <= 5'd23/*23:xpc10:23*/;
                       TSPte2_13_V_0 <= 33'h1ffffffff&32'd0;
                       phase <= 33'h1ffffffff&32'd8+32'd256*TSPru0_12_V_1;
                       end 
                      
              5'd23/*23:US*/: if ((TSPte2_13_V_0<2'd2))  begin 
                       xpc10 <= 5'd30/*30:xpc10:30*/;
                       TSPte2_13_V_2 <= 33'h1ffffffff&32'd0;
                       TSPte2_13_V_1 <= 33'h1ffffffff&((TSPru0_12_V_1+TSPte2_13_V_0)%2'd2);
                       end 
                       else  begin 
                       xpc10 <= 5'd24/*24:xpc10:24*/;
                       A_UINT_CC_SCALbx36_crc_reg <= 33'h1ffffffff&-32'd1;
                       phase <= 33'h1ffffffff&32'd10+32'd256*TSPru0_12_V_1;
                       end 
                      
              5'd25/*25:US*/:  begin 
                  if ((TSPcr2_16_V_1>=(33'h1ffffffff&32'h4d))) $display("step %d crc is %d", TSPru0_12_V_1, A_UINT_CC_SCALbx36_crc_reg
                      );
                       else $display("process unit word %d word=%d", A_UINT_CC_SCALbx36_byteno, 33'h1ffffffff&A_64_SS_CC_SCALbx54_ARB0
                      [(65'h1ffffffffffffffff&TSPcr2_16_V_1)+(65'h1ffffffffffffffff&TSPcr2_16_V_0)*A_SINT_CC_SCALbx42_d2dim0]);
                  if ((TSPcr2_16_V_1<(33'h1ffffffff&32'h4d)))  begin 
                           xpc10 <= 5'd26/*26:xpc10:26*/;
                           A_UINT_CC_SCALbx36_byteno <= 33'h1ffffffff&32'd1+A_UINT_CC_SCALbx36_byteno;
                           TCpr0_13_V_0 <= 9'h1ff&8'd255&(A_UINT_CC_SCALbx36_crc_reg>>5'd24);
                           TSPcr2_16_V_2 <= 65'h1ffffffffffffffff&A_64_SS_CC_SCALbx54_ARB0[(65'h1ffffffffffffffff&TSPcr2_16_V_1)+(65'h1ffffffffffffffff
                          &TSPcr2_16_V_0)*A_SINT_CC_SCALbx42_d2dim0];

                           end 
                           else  begin 
                           xpc10 <= 5'd19/*19:xpc10:19*/;
                           TSPru0_12_V_1 <= 33'h1ffffffff&32'd1+TSPru0_12_V_1;
                           d_monitor <= 65'h1ffffffffffffffff&A_UINT_CC_SCALbx36_crc_reg;
                           end 
                           end 
                  
              5'd31/*31:US*/:  begin 
                  $write("%d %d : %d   ", TSPte2_13_V_1, TSPte2_13_V_2, 65'h1ffffffffffffffff&A_64_SS_CC_SCALbx54_ARB0[(65'h1ffffffffffffffff
                  &TSPte2_13_V_2)+(65'h1ffffffffffffffff&TSPte2_13_V_1)*A_SINT_CC_SCALbx42_d2dim0]);
                  $display("");
                   end 
                  
              6'd32/*32:US*/: if (((65'h1ffffffffffffffff&(33'h1ffffffff&-32'd2)+A_64_SS_CC_SCALbx58_ARD0[(65'h1ffffffffffffffff&64'd1
              +TSPne2_10_V_3)+(65'h1ffffffffffffffff&TSPne2_10_V_0)*A_SINT_CC_SCALbx46_d2dim0])<A_64_SS_CC_SCALbx52_ARA0[(65'h1ffffffffffffffff
              &64'd1+TSPne2_10_V_3)+(65'h1ffffffffffffffff&TSPne2_10_V_0)*A_SINT_CC_SCALbx40_d2dim0]))  begin 
                       xpc10 <= 6'd33/*33:xpc10:33*/;
                       TSPne2_10_V_4 <= 33'h1ffffffff&A_SINT_CC_SCALbx26_ARJ0[TSPne2_10_V_3];
                       A_64_SS_CC_SCALbx58_ARD0[(65'h1ffffffffffffffff&64'd1+TSPne2_10_V_3)+(65'h1ffffffffffffffff&TSPne2_10_V_1)*A_SINT_CC_SCALbx46_d2dim0
                      ] <= 65'h1ffffffffffffffff&A_64_SS_CC_SCALbx52_ARA0[(65'h1ffffffffffffffff&64'd1+TSPne2_10_V_3)+(65'h1ffffffffffffffff
                      &TSPne2_10_V_0)*A_SINT_CC_SCALbx40_d2dim0];

                       end 
                       else  begin 
                       xpc10 <= 6'd33/*33:xpc10:33*/;
                       TSPne2_10_V_4 <= 33'h1ffffffff&A_SINT_CC_SCALbx26_ARJ0[TSPne2_10_V_3];
                       A_64_SS_CC_SCALbx58_ARD0[(65'h1ffffffffffffffff&64'd1+TSPne2_10_V_3)+(65'h1ffffffffffffffff&TSPne2_10_V_1)*A_SINT_CC_SCALbx46_d2dim0
                      ] <= 65'h1ffffffffffffffff&(33'h1ffffffff&-32'd2)+A_64_SS_CC_SCALbx58_ARD0[(65'h1ffffffffffffffff&64'd1+TSPne2_10_V_3
                      )+(65'h1ffffffffffffffff&TSPne2_10_V_0)*A_SINT_CC_SCALbx46_d2dim0];

                       end 
                      
              6'd39/*39:US*/:  begin 
                   xpc10 <= 5'd18/*18:xpc10:18*/;
                   TSPsw1_2_V_1 <= 33'h1ffffffff&32'd1+TSPsw1_2_V_1;
                   A_64_SS_CC_SCALbx52_ARA0[(65'h1ffffffffffffffff&TSPsw1_2_V_1)+(33'h1ffffffff&32'd0)*A_SINT_CC_SCALbx40_d2dim0] <= 65'h1ffffffffffffffff
                  &-64'd10;

                   A_64_SS_CC_SCALbx54_ARB0[(65'h1ffffffffffffffff&TSPsw1_2_V_1)+(33'h1ffffffff&32'd0)*A_SINT_CC_SCALbx42_d2dim0] <= 33'h1ffffffff
                  &32'd0;

                   A_64_SS_CC_SCALbx56_ARC0[(65'h1ffffffffffffffff&TSPsw1_2_V_1)+(33'h1ffffffff&32'd0)*A_SINT_CC_SCALbx44_d2dim0] <= 33'h1ffffffff
                  &32'd0;

                   A_64_SS_CC_SCALbx58_ARD0[(65'h1ffffffffffffffff&TSPsw1_2_V_1)+(33'h1ffffffff&32'd0)*A_SINT_CC_SCALbx46_d2dim0] <= 33'h1ffffffff
                  &32'd0;

                   end 
                  
              6'd40/*40:US*/:  begin 
                   xpc10 <= 5'd17/*17:xpc10:17*/;
                   TSPsw1_2_V_0 <= 33'h1ffffffff&32'd1+TSPsw1_2_V_0;
                   d_monitor <= 65'h1ffffffffffffffff&TSPsw1_2_V_0;
                   A_64_SS_CC_SCALbx52_ARA0[(33'h1ffffffff&32'd0)+(65'h1ffffffffffffffff&TSPsw1_2_V_0)*A_SINT_CC_SCALbx40_d2dim0] <= 65'h1ffffffffffffffff
                  &-64'd10;

                   A_64_SS_CC_SCALbx54_ARB0[(33'h1ffffffff&32'd0)+(65'h1ffffffffffffffff&TSPsw1_2_V_0)*A_SINT_CC_SCALbx42_d2dim0] <= 33'h1ffffffff
                  &32'd0;

                   A_64_SS_CC_SCALbx56_ARC0[(33'h1ffffffff&32'd0)+(65'h1ffffffffffffffff&TSPsw1_2_V_0)*A_SINT_CC_SCALbx44_d2dim0] <= 33'h1ffffffff
                  &32'd0;

                   A_64_SS_CC_SCALbx58_ARD0[(33'h1ffffffff&32'd0)+(65'h1ffffffffffffffff&TSPsw1_2_V_0)*A_SINT_CC_SCALbx46_d2dim0] <= 33'h1ffffffff
                  &32'd0;

                   end 
                  endcase
              if ((A_16_SS_CC_SCALbx10_ARA0[TSPru0_12_V_1]==A_16_SS_CC_SCALbx12_ARB0[TSPen0_17_V_0]))  begin if ((xpc10==6'd38/*38:US*/)) 
                           begin 
                           xpc10 <= 5'd21/*21:xpc10:21*/;
                           TSPe0_SPILL_256 <= 33'h1ffffffff&TSPen0_17_V_0;
                           end 
                           end 
                   else if ((xpc10==6'd38/*38:US*/))  begin 
                           xpc10 <= 5'd20/*20:xpc10:20*/;
                           TSPen0_17_V_0 <= 33'h1ffffffff&32'd1+TSPen0_17_V_0;
                           end 
                          
              case (xpc10)

              5'd26/*26:US*/:  begin 
                   xpc10 <= 5'd27/*27:xpc10:27*/;
                   A_UINT_CC_SCALbx36_byteno <= 33'h1ffffffff&32'd1+A_UINT_CC_SCALbx36_byteno;
                   TCpr0_21_V_0 <= 9'h1ff&8'd255&((33'h1ffffffff&-32'd1&A_UINT_CC_SCALbx34_ARA0[9'h1ff&8'd255&33'h1ffffffff&TSPcr2_16_V_2
                  ]^A_UINT_CC_SCALbx34_ARA0[TCpr0_13_V_0]^{A_UINT_CC_SCALbx36_crc_reg, 8'd0})>>5'd24);

                   A_UINT_CC_SCALbx36_crc_reg <= 33'h1ffffffff&-32'd1&A_UINT_CC_SCALbx34_ARA0[9'h1ff&8'd255&33'h1ffffffff&TSPcr2_16_V_2
                  ]^A_UINT_CC_SCALbx34_ARA0[TCpr0_13_V_0]^{A_UINT_CC_SCALbx36_crc_reg, 8'd0};

                   end 
                  
              5'd27/*27:US*/:  begin 
                   xpc10 <= 5'd28/*28:xpc10:28*/;
                   A_UINT_CC_SCALbx36_byteno <= 33'h1ffffffff&32'd1+A_UINT_CC_SCALbx36_byteno;
                   TCpr0_29_V_0 <= 9'h1ff&8'd255&((33'h1ffffffff&-32'd1&A_UINT_CC_SCALbx34_ARA0[9'h1ff&8'd255&((33'h1ffffffff&TSPcr2_16_V_2
                  )>>4'd8)]^A_UINT_CC_SCALbx34_ARA0[TCpr0_21_V_0]^{A_UINT_CC_SCALbx36_crc_reg, 8'd0})>>5'd24);

                   A_UINT_CC_SCALbx36_crc_reg <= 33'h1ffffffff&-32'd1&A_UINT_CC_SCALbx34_ARA0[9'h1ff&8'd255&((33'h1ffffffff&TSPcr2_16_V_2
                  )>>4'd8)]^A_UINT_CC_SCALbx34_ARA0[TCpr0_21_V_0]^{A_UINT_CC_SCALbx36_crc_reg, 8'd0};

                   end 
                  
              5'd28/*28:US*/:  begin 
                   xpc10 <= 5'd29/*29:xpc10:29*/;
                   A_UINT_CC_SCALbx36_byteno <= 33'h1ffffffff&32'd1+A_UINT_CC_SCALbx36_byteno;
                   TCpr0_35_V_0 <= 9'h1ff&8'd255&((33'h1ffffffff&-32'd1&A_UINT_CC_SCALbx34_ARA0[9'h1ff&8'd255&((33'h1ffffffff&TSPcr2_16_V_2
                  )>>5'd16)]^A_UINT_CC_SCALbx34_ARA0[TCpr0_29_V_0]^{A_UINT_CC_SCALbx36_crc_reg, 8'd0})>>5'd24);

                   A_UINT_CC_SCALbx36_crc_reg <= 33'h1ffffffff&-32'd1&A_UINT_CC_SCALbx34_ARA0[9'h1ff&8'd255&((33'h1ffffffff&TSPcr2_16_V_2
                  )>>5'd16)]^A_UINT_CC_SCALbx34_ARA0[TCpr0_29_V_0]^{A_UINT_CC_SCALbx36_crc_reg, 8'd0};

                   end 
                  
              5'd31/*31:US*/:  begin 
                   xpc10 <= 5'd30/*30:xpc10:30*/;
                   TSPte2_13_V_2 <= 33'h1ffffffff&32'd1+TSPte2_13_V_2;
                   end 
                  
              6'd33/*33:US*/: if (((65'h1ffffffffffffffff&(33'h1ffffffff&-32'd2)+A_64_SS_CC_SCALbx56_ARC0[(65'h1ffffffffffffffff&TSPne2_10_V_3
              )+(65'h1ffffffffffffffff&TSPne2_10_V_1)*A_SINT_CC_SCALbx44_d2dim0])<A_64_SS_CC_SCALbx52_ARA0[(65'h1ffffffffffffffff&TSPne2_10_V_3
              )+(65'h1ffffffffffffffff&TSPne2_10_V_1)*A_SINT_CC_SCALbx40_d2dim0]))  begin 
                       xpc10 <= 6'd34/*34:xpc10:34*/;
                       A_64_SS_CC_SCALbx56_ARC0[(65'h1ffffffffffffffff&64'd1+TSPne2_10_V_3)+(65'h1ffffffffffffffff&TSPne2_10_V_1)*A_SINT_CC_SCALbx44_d2dim0
                      ] <= 65'h1ffffffffffffffff&A_64_SS_CC_SCALbx52_ARA0[(65'h1ffffffffffffffff&TSPne2_10_V_3)+(65'h1ffffffffffffffff
                      &TSPne2_10_V_1)*A_SINT_CC_SCALbx40_d2dim0];

                       end 
                       else  begin 
                       xpc10 <= 6'd34/*34:xpc10:34*/;
                       A_64_SS_CC_SCALbx58_ARD0[(65'h1ffffffffffffffff&64'd1+TSPne2_10_V_3)+(65'h1ffffffffffffffff&TSPne2_10_V_1)*A_SINT_CC_SCALbx46_d2dim0
                      ] <= 65'h1ffffffffffffffff&(33'h1ffffffff&-32'd2)+A_64_SS_CC_SCALbx56_ARC0[(65'h1ffffffffffffffff&TSPne2_10_V_3
                      )+(65'h1ffffffffffffffff&TSPne2_10_V_1)*A_SINT_CC_SCALbx44_d2dim0];

                       end 
                      
              6'd34/*34:US*/: if ((A_64_SS_CC_SCALbx56_ARC0[(65'h1ffffffffffffffff&TSPne2_10_V_3)+(65'h1ffffffffffffffff&TSPne2_10_V_0
              )*A_SINT_CC_SCALbx44_d2dim0]<A_64_SS_CC_SCALbx58_ARD0[(65'h1ffffffffffffffff&TSPne2_10_V_3)+(65'h1ffffffffffffffff&TSPne2_10_V_0
              )*A_SINT_CC_SCALbx46_d2dim0]))  begin 
                       xpc10 <= 6'd35/*35:xpc10:35*/;
                       TSPne2_10_V_7 <= 65'h1ffffffffffffffff&A_64_SS_CC_SCALbx58_ARD0[(65'h1ffffffffffffffff&TSPne2_10_V_3)+(65'h1ffffffffffffffff
                      &TSPne2_10_V_0)*A_SINT_CC_SCALbx46_d2dim0];

                       end 
                       else  begin 
                       xpc10 <= 6'd35/*35:xpc10:35*/;
                       TSPne2_10_V_7 <= 65'h1ffffffffffffffff&A_64_SS_CC_SCALbx56_ARC0[(65'h1ffffffffffffffff&TSPne2_10_V_3)+(65'h1ffffffffffffffff
                      &TSPne2_10_V_0)*A_SINT_CC_SCALbx44_d2dim0];

                       end 
                      
              6'd36/*36:US*/: if (((65'h1ffffffffffffffff&TSPne2_10_V_7+A_SINT_CC_SCALbx16_ARA0[(65'h1ffffffffffffffff&TSPne2_10_V_2)+
              (65'h1ffffffffffffffff&TSPne2_10_V_4)*A_SINT_CC_SCALbx32_d2dim0])<(33'h1ffffffff&32'd0)))  begin 
                       xpc10 <= 6'd37/*37:xpc10:37*/;
                       A_64_SS_CC_SCALbx54_ARB0[(65'h1ffffffffffffffff&64'd1+TSPne2_10_V_3)+(65'h1ffffffffffffffff&TSPne2_10_V_1)*A_SINT_CC_SCALbx42_d2dim0
                      ] <= 33'h1ffffffff&32'd0;

                       end 
                       else  begin 
                       xpc10 <= 6'd37/*37:xpc10:37*/;
                       A_64_SS_CC_SCALbx54_ARB0[(65'h1ffffffffffffffff&64'd1+TSPne2_10_V_3)+(65'h1ffffffffffffffff&TSPne2_10_V_1)*A_SINT_CC_SCALbx42_d2dim0
                      ] <= 65'h1ffffffffffffffff&TSPne2_10_V_7+A_SINT_CC_SCALbx16_ARA0[(65'h1ffffffffffffffff&TSPne2_10_V_2)+(65'h1ffffffffffffffff
                      &TSPne2_10_V_4)*A_SINT_CC_SCALbx32_d2dim0];

                       end 
                      endcase
              if ((A_16_SS_CC_SCALbx12_ARB0[TSPen1_8_V_0]==A_16_SS_CC_SCALbx14_ARC0[TSPin0_6_V_0]))  begin if ((xpc10==2'd2/*2:US*/)) 
                           begin 
                           xpc10 <= 2'd3/*3:xpc10:3*/;
                           TSPe1_SPILL_256 <= 33'h1ffffffff&TSPen1_8_V_0;
                           end 
                           end 
                   else if ((xpc10==2'd2/*2:US*/))  begin 
                           xpc10 <= 6'd41/*41:xpc10:41*/;
                           TSPen1_8_V_0 <= 33'h1ffffffff&32'd1+TSPen1_8_V_0;
                           end 
                          
              case (xpc10)

              3'd6/*6:US*/:  begin 
                   xpc10 <= 3'd7/*7:xpc10:7*/;
                   A_UINT_CC_SCALbx38_crc_reg <= 33'h1ffffffff&-32'd1;
                   end 
                  
              3'd7/*7:US*/:  xpc10 <= 4'd8/*8:xpc10:8*/;

              4'd8/*8:US*/:  xpc10 <= 4'd9/*9:xpc10:9*/;

              4'd9/*9:US*/:  xpc10 <= 4'd10/*10:xpc10:10*/;

              4'd10/*10:US*/:  begin 
                   xpc10 <= 4'd11/*11:xpc10:11*/;
                   A_UINT_CC_SCALbx38_crc_reg <= 33'h1ffffffff&-32'd1&A_UINT_CC_SCALbx34_ARA0[32'd255]^A_UINT_CC_SCALbx34_ARA0[32'd1]
                  ^{A_UINT_CC_SCALbx38_crc_reg, 8'd0};

                   end 
                  
              4'd11/*11:US*/:  begin 
                   xpc10 <= 4'd12/*12:xpc10:12*/;
                   TCpr0_40_V_0 <= 9'h1ff&8'd255&(A_UINT_CC_SCALbx38_crc_reg>>5'd24);
                   end 
                  
              4'd12/*12:US*/:  begin 
                   xpc10 <= 4'd13/*13:xpc10:13*/;
                   A_UINT_CC_SCALbx38_crc_reg <= 33'h1ffffffff&-32'd1&A_UINT_CC_SCALbx34_ARA0[32'd128]^A_UINT_CC_SCALbx34_ARA0[TCpr0_40_V_0
                  ]^{A_UINT_CC_SCALbx38_crc_reg, 8'd0};

                   end 
                  
              4'd13/*13:US*/:  begin 
                   xpc10 <= 4'd14/*14:xpc10:14*/;
                   TCpr0_44_V_0 <= 9'h1ff&8'd255&(A_UINT_CC_SCALbx38_crc_reg>>5'd24);
                   end 
                  
              4'd14/*14:US*/:  begin 
                   xpc10 <= 4'd15/*15:xpc10:15*/;
                   A_UINT_CC_SCALbx38_crc_reg <= 33'h1ffffffff&-32'd1&A_UINT_CC_SCALbx34_ARA0[32'd1]^A_UINT_CC_SCALbx34_ARA0[TCpr0_44_V_0
                  ]^{A_UINT_CC_SCALbx38_crc_reg, 8'd0};

                   end 
                  
              5'd16/*16:US*/:  begin 
                   xpc10 <= 5'd17/*17:xpc10:17*/;
                   TSPsw1_2_V_0 <= 33'h1ffffffff&32'd0;
                   end 
                  
              5'd17/*17:US*/: if ((TSPsw1_2_V_0<2'd2))  xpc10 <= 6'd40/*40:xpc10:40*/;
                   else  begin 
                       xpc10 <= 5'd18/*18:xpc10:18*/;
                       TSPsw1_2_V_1 <= 33'h1ffffffff&32'd1;
                       end 
                      
              5'd18/*18:US*/: if ((TSPsw1_2_V_1<7'd78))  xpc10 <= 6'd39/*39:xpc10:39*/;
                   else  begin 
                       xpc10 <= 5'd19/*19:xpc10:19*/;
                       TSPru0_12_V_1 <= 33'h1ffffffff&32'd0;
                       end 
                      
              5'd20/*20:US*/: if ((TSPen0_17_V_0<5'd20))  xpc10 <= 6'd38/*38:xpc10:38*/;
                   else  begin 
                       xpc10 <= 5'd21/*21:xpc10:21*/;
                       TSPe0_SPILL_256 <= 33'h1ffffffff&32'd0;
                       end 
                      
              5'd21/*21:US*/:  begin 
                   xpc10 <= 5'd22/*22:xpc10:22*/;
                   TSPne2_10_V_3 <= 33'h1ffffffff&32'd0;
                   TSPne2_10_V_2 <= 33'h1ffffffff&TSPe0_SPILL_256;
                   end 
                  
              5'd24/*24:US*/:  begin 
                   xpc10 <= 5'd25/*25:xpc10:25*/;
                   TSPcr2_16_V_1 <= 33'h1ffffffff&32'd0;
                   TSPcr2_16_V_0 <= 33'h1ffffffff&((32'd1+TSPru0_12_V_1)%2'd2);
                   end 
                  
              5'd29/*29:US*/:  begin 
                   xpc10 <= 5'd25/*25:xpc10:25*/;
                   TSPcr2_16_V_1 <= 33'h1ffffffff&32'd1+TSPcr2_16_V_1;
                   A_UINT_CC_SCALbx36_crc_reg <= 33'h1ffffffff&-32'd1&A_UINT_CC_SCALbx34_ARA0[9'h1ff&8'd255&33'h1ffffffff&TSPcr2_16_V_2
                  ]^A_UINT_CC_SCALbx34_ARA0[TCpr0_35_V_0]^{A_UINT_CC_SCALbx36_crc_reg, 8'd0};

                   end 
                  
              5'd30/*30:US*/: if ((TSPte2_13_V_2<(33'h1ffffffff&32'h4d)))  xpc10 <= 5'd31/*31:xpc10:31*/;
                   else  begin 
                       xpc10 <= 5'd23/*23:xpc10:23*/;
                       TSPte2_13_V_0 <= 33'h1ffffffff&32'd1+TSPte2_13_V_0;
                       end 
                      
              6'd35/*35:US*/: if ((TSPne2_10_V_7<A_64_SS_CC_SCALbx54_ARB0[(65'h1ffffffffffffffff&TSPne2_10_V_3)+(65'h1ffffffffffffffff
              &TSPne2_10_V_0)*A_SINT_CC_SCALbx42_d2dim0]))  begin 
                       xpc10 <= 6'd36/*36:xpc10:36*/;
                       TSPne2_10_V_7 <= 65'h1ffffffffffffffff&A_64_SS_CC_SCALbx54_ARB0[(65'h1ffffffffffffffff&TSPne2_10_V_3)+(65'h1ffffffffffffffff
                      &TSPne2_10_V_0)*A_SINT_CC_SCALbx42_d2dim0];

                       end 
                       else  xpc10 <= 6'd36/*36:xpc10:36*/;

              6'd37/*37:US*/:  begin 
                   xpc10 <= 5'd22/*22:xpc10:22*/;
                   TSPne2_10_V_3 <= 33'h1ffffffff&64'd1+TSPne2_10_V_3;
                   A_64_SS_CC_SCALbx52_ARA0[(65'h1ffffffffffffffff&64'd1+TSPne2_10_V_3)+(65'h1ffffffffffffffff&TSPne2_10_V_1)*A_SINT_CC_SCALbx40_d2dim0
                  ] <= 65'h1ffffffffffffffff&(65'h1ffffffffffffffff&-64'd10)+A_64_SS_CC_SCALbx54_ARB0[(65'h1ffffffffffffffff&64'd1+TSPne2_10_V_3
                  )+(65'h1ffffffffffffffff&TSPne2_10_V_1)*A_SINT_CC_SCALbx42_d2dim0];

                   end 
                  
              6'd41/*41:US*/: if ((TSPen1_8_V_0<5'd20))  xpc10 <= 1'd1/*1:xpc10:1*/;
                   else  begin 
                       xpc10 <= 2'd3/*3:xpc10:3*/;
                       TSPe1_SPILL_256 <= 33'h1ffffffff&32'd0;
                       end 
                      endcase
              if ((xpc10==1'd1/*1:US*/))  xpc10 <= 2'd2/*2:xpc10:2*/;
                  if ((xpc10==3'd5/*5:US*/))  xpc10 <= 3'd6/*6:xpc10:6*/;
                   end 
              //End structure HPR sw_test.exe


       end 
      

//Total area 0
// 1 vectors of width 6
// 8 vectors of width 32
// 6 vectors of width 8
// 2 vectors of width 64
// 338 array locations of width 16
// 1385 array locations of width 32
// 624 array locations of width 64
// 608 bits in scalar variables
// Total state bits in module = 90710 bits.
// Total number of leaf cells = 0
endmodule

//  
// LCP delay estimations included: turn off with -vnl-lcp-delay-estimate=disable
// eof (HPR L/S Verilog)
