

// CBG Orangepath HPR L/S System

// Verilog output file generated at 25/09/2016 22:38:42
// Kiwi Scientific Acceleration (KiwiC .net/CIL/C# to Verilog/SystemC compiler): Version alpha 0.2.16f : 22nd-September-2016 Linux/X86_64:koo
//  /home/djg11/d320/hprls/kiwipro/kiwic/distro/lib/kiwic.exe -vnl-resets=synchronous -restructure2=disable -vnl-roundtrip=disable -kiwic-cil-dump=combined -kiwic-kcode-dump=enable -bevelab-default-pause-mode=soft -bevelab-soft-pause-threshold=10 dfsin.exe -vnl=dfsin.v -vnl-resets=synchronous ../softfloat.dll
`timescale 1ns/1ns


module dfsin(output reg done, input [31:0] dfsin_arg, output [31:0] dfsin_result, input clk, input reset);
function signed [15:0] rtl_signed_bitextract9;
   input [63:0] arg;
   rtl_signed_bitextract9 = $signed(arg[15:0]);
   endfunction

function signed [15:0] rtl_signed_bitextract0;
   input [31:0] arg;
   rtl_signed_bitextract0 = $signed(arg[15:0]);
   endfunction

function  rtl_unsigned_bitextract8;
   input [31:0] arg;
   rtl_unsigned_bitextract8 = $unsigned(arg[0:0]);
   endfunction

function  rtl_unsigned_bitextract5;
   input [31:0] arg;
   rtl_unsigned_bitextract5 = $unsigned(arg[0:0]);
   endfunction

function [7:0] rtl_unsigned_bitextract3;
   input [31:0] arg;
   rtl_unsigned_bitextract3 = $unsigned(arg[7:0]);
   endfunction

function [31:0] rtl_unsigned_bitextract1;
   input [63:0] arg;
   rtl_unsigned_bitextract1 = $unsigned(arg[31:0]);
   endfunction

function signed [63:0] rtl_sign_extend11;
   input [15:0] arg;
   rtl_sign_extend11 = { {48{arg[15]}}, arg[15:0] };
   endfunction

function signed [31:0] rtl_sign_extend10;
   input [7:0] arg;
   rtl_sign_extend10 = { {24{arg[7]}}, arg[7:0] };
   endfunction

function signed [31:0] rtl_sign_extend6;
   input argbit;
   rtl_sign_extend6 = { {32{argbit}} };
   endfunction

function signed [63:0] rtl_sign_extend4;
   input [31:0] arg;
   rtl_sign_extend4 = { {32{arg[31]}}, arg[31:0] };
   endfunction

function signed [31:0] rtl_sign_extend2;
   input [15:0] arg;
   rtl_sign_extend2 = { {16{arg[15]}}, arg[15:0] };
   endfunction

function [63:0] rtl_unsigned_extend7;
   input [31:0] arg;
   rtl_unsigned_extend7 = { 32'b0, arg[31:0] };
   endfunction

  integer dfsin_gloops;
  integer Tdbm0_3_V_0;
  integer Tdbm0_3_V_1;
  reg [63:0] Tdsi3_5_V_0;
  reg [63:0] Tdsi3_5_V_1;
  integer Tdsi3_5_V_2;
  reg [63:0] Tsfl0_9_V_8;
  reg [63:0] Tsfl0_9_V_9;
  reg [63:0] Tsfl0_9_V_6;
  reg signed [15:0] Tsfl0_9_V_3;
  reg Tsfl0_9_V_0;
  reg [63:0] Tsfl0_9_V_7;
  reg signed [15:0] Tsfl0_9_V_4;
  reg Tsfl0_9_V_1;
  reg Tsfl0_9_V_2;
  reg [63:0] Tsf0_SPILL_256;
  reg [63:0] Tspr4_3_V_0;
  reg [63:0] Tspr4_3_V_1;
  integer Tsf0SPILL10_256;
  reg Tspr4_3_V_2;
  reg Tspr4_3_V_3;
  integer Tsf0SPILL12_256;
  reg Tspr4_3_V_4;
  reg [63:0] Tspr11_2_V_0;
  reg [63:0] Tspr11_2_V_1;
  reg Tspr11_2_V_2;
  reg Tspr11_2_V_3;
  reg Tspr11_2_V_4;
  reg [63:0] Tsco0_2_V_0;
  reg [7:0] Tsco0_2_V_1;
  reg [31:0] Tsco3_7_V_0;
  reg [7:0] Tsco3_7_V_1;
  integer Tsno19_4_V_0;
  integer Tsno23_4_V_0;
  reg signed [15:0] Tsfl0_9_V_5;
  reg [31:0] Tsmu24_24_V_1;
  reg [31:0] Tsmu24_24_V_0;
  reg [31:0] Tsmu24_24_V_3;
  reg [31:0] Tsmu24_24_V_2;
  reg [63:0] Tsmu24_24_V_7;
  reg [63:0] Tsmu24_24_V_5;
  reg [63:0] Tsmu24_24_V_6;
  reg [63:0] Tsmu24_24_V_4;
  reg [63:0] fastspilldup16;
  reg [63:0] Tsm24_SPILL_264;
  reg [63:0] Tsm24_SPILL_257;
  reg signed [63:0] Tsm24_SPILL_259;
  reg [63:0] fastspilldup18;
  reg [63:0] Tsm24_SPILL_263;
  reg [63:0] Tsm24_SPILL_260;
  reg signed [63:0] Tsm24_SPILL_262;
  reg [63:0] fastspilldup20;
  reg [63:0] Tsf0_SPILL_260;
  reg [63:0] Tsf0_SPILL_257;
  reg signed [63:0] Tsf0_SPILL_259;
  reg signed [15:0] Tsro29_4_V_0;
  reg [63:0] Tsro29_4_V_1;
  reg signed [15:0] Tsro29_4_V_5;
  reg signed [15:0] Tsro29_4_V_6;
  reg [63:0] Tssh18_7_V_0;
  reg [63:0] fastspilldup24;
  reg [63:0] Tss18_SPILL_259;
  reg [63:0] Tss18_SPILL_256;
  reg signed [63:0] Tss18_SPILL_258;
  reg [63:0] Tss18_SPILL_257;
  reg signed [63:0] Tss18_SPILL_260;
  reg [63:0] fastspilldup22;
  reg [63:0] Tsr29_SPILL_260;
  reg [63:0] Tsr29_SPILL_256;
  reg signed [63:0] Tsr29_SPILL_258;
  reg [63:0] Tsr29_SPILL_257;
  reg [63:0] Tsr29_SPILL_259;
  reg signed [63:0] Tsp27_SPILL_256;
  reg [63:0] Tsfl0_10_V_0;
  reg [63:0] Tdsi3_5_V_3;
  reg [63:0] Tsfl1_7_V_8;
  reg [63:0] Tsfl1_7_V_9;
  reg [63:0] Tsfl1_7_V_6;
  reg signed [15:0] Tsfl1_7_V_3;
  reg Tsfl1_7_V_0;
  reg [63:0] Tsfl1_7_V_7;
  reg signed [15:0] Tsfl1_7_V_4;
  reg Tsfl1_7_V_1;
  reg Tsfl1_7_V_2;
  reg [63:0] Tsf1_SPILL_256;
  reg signed [15:0] Tsfl1_7_V_5;
  reg [63:0] fastspilldup26;
  reg [63:0] fastspilldup28;
  reg [63:0] fastspilldup30;
  reg [63:0] Tsf1_SPILL_260;
  reg [63:0] Tsf1_SPILL_257;
  reg signed [63:0] Tsf1_SPILL_259;
  reg [63:0] fastspilldup34;
  reg [63:0] fastspilldup32;
  reg [63:0] Tsi1_SPILL_256;
  reg Tsin1_17_V_0;
  integer Tsi1_SPILL_257;
  reg [31:0] Tsin1_17_V_1;
  reg [31:0] Tsco5_4_V_0;
  reg [7:0] Tsco5_4_V_1;
  integer Tsin1_17_V_3;
  reg [63:0] Tsin1_17_V_2;
  reg signed [63:0] Tsp5_SPILL_256;
  reg [63:0] Tsfl1_18_V_6;
  reg signed [15:0] Tsfl1_18_V_3;
  reg Tsfl1_18_V_0;
  reg [63:0] Tsfl1_18_V_7;
  reg signed [15:0] Tsfl1_18_V_4;
  reg Tsfl1_18_V_1;
  reg Tsfl1_18_V_2;
  reg [63:0] Tspr2_2_V_0;
  reg [63:0] Tspr2_2_V_1;
  reg Tspr2_2_V_2;
  reg Tspr2_2_V_3;
  reg Tspr2_2_V_4;
  reg [63:0] Tsf1SPILL10_256;
  reg [63:0] Tspr5_2_V_0;
  reg [63:0] Tspr5_2_V_1;
  reg Tspr5_2_V_2;
  reg Tspr5_2_V_3;
  reg Tspr5_2_V_4;
  reg [63:0] Tspr10_2_V_0;
  reg [63:0] Tspr10_2_V_1;
  reg Tspr10_2_V_2;
  reg Tspr10_2_V_3;
  reg Tspr10_2_V_4;
  integer Tsno18_4_V_0;
  integer Tsno22_4_V_0;
  reg signed [15:0] Tsfl1_18_V_5;
  reg [63:0] Tses25_5_V_0;
  reg [63:0] Tse25_SPILL_257;
  reg [63:0] Tses25_5_V_6;
  reg [31:0] Tsmu5_7_V_1;
  reg [31:0] Tsmu5_7_V_0;
  reg [31:0] Tsmu5_7_V_3;
  reg [31:0] Tsmu5_7_V_2;
  reg [63:0] Tsmu5_7_V_7;
  reg [63:0] Tsmu5_7_V_5;
  reg [63:0] Tsmu5_7_V_6;
  reg [63:0] Tsmu5_7_V_4;
  reg [63:0] fastspilldup36;
  reg [63:0] Tsm5_SPILL_264;
  reg [63:0] Tsm5_SPILL_257;
  reg signed [63:0] Tsm5_SPILL_259;
  reg [63:0] fastspilldup38;
  reg [63:0] Tsm5_SPILL_263;
  reg [63:0] Tsm5_SPILL_260;
  reg signed [63:0] Tsm5_SPILL_262;
  reg [63:0] Tses25_5_V_5;
  reg [63:0] Tses25_5_V_4;
  reg [63:0] Tses25_5_V_3;
  reg [63:0] fastspilldup40;
  reg [63:0] Tss5_SPILL_262;
  reg [63:0] Tss5_SPILL_257;
  reg signed [63:0] Tss5_SPILL_260;
  reg [63:0] Tss5_SPILL_259;
  reg [63:0] Tses25_5_V_2;
  reg [63:0] fastspilldup44;
  reg [63:0] Tse25_SPILL_261;
  reg [63:0] Tse25_SPILL_258;
  reg [63:0] Tse25_SPILL_260;
  reg [63:0] Tsfl1_18_V_8;
  reg [31:0] Tsmu26_4_V_1;
  reg [31:0] Tsmu26_4_V_0;
  reg [31:0] Tsmu26_4_V_3;
  reg [31:0] Tsmu26_4_V_2;
  reg [63:0] Tsmu26_4_V_7;
  reg [63:0] Tsmu26_4_V_5;
  reg [63:0] Tsmu26_4_V_6;
  reg [63:0] Tsmu26_4_V_4;
  reg [63:0] fastspilldup46;
  reg [63:0] Tsm26_SPILL_264;
  reg [63:0] Tsm26_SPILL_257;
  reg signed [63:0] Tsm26_SPILL_259;
  reg [63:0] fastspilldup48;
  reg [63:0] Tsm26_SPILL_263;
  reg [63:0] Tsm26_SPILL_260;
  reg signed [63:0] Tsm26_SPILL_262;
  reg [63:0] Tsfl1_18_V_12;
  reg [63:0] Tsfl1_18_V_11;
  reg [63:0] Tsfl1_18_V_10;
  reg [63:0] fastspilldup50;
  reg [63:0] Tss26_SPILL_262;
  reg [63:0] Tss26_SPILL_257;
  reg signed [63:0] Tss26_SPILL_260;
  reg [63:0] Tss26_SPILL_259;
  reg [63:0] Tsfl1_18_V_9;
  reg [63:0] fastspilldup54;
  reg [63:0] Tsf1SPILL10_260;
  reg [63:0] Tsf1SPILL10_257;
  reg signed [63:0] Tsf1SPILL10_259;
  reg [63:0] Tsad27_13_V_0;
  reg [63:0] fastspilldup52;
  reg [63:0] Tsa27_SPILL_262;
  reg [63:0] Tsa27_SPILL_257;
  reg signed [63:0] Tsa27_SPILL_260;
  reg [63:0] Tsa27_SPILL_259;
  reg signed [15:0] Tsro33_4_V_0;
  reg [63:0] Tsro33_4_V_1;
  reg signed [15:0] Tsro33_4_V_5;
  reg signed [15:0] Tsro33_4_V_6;
  reg [63:0] fastspilldup58;
  reg [63:0] fastspilldup56;
  reg [63:0] Tsr33_SPILL_260;
  reg [63:0] Tsr33_SPILL_256;
  reg signed [63:0] Tsr33_SPILL_258;
  reg [63:0] Tsr33_SPILL_257;
  reg [63:0] Tsr33_SPILL_259;
  integer Tse0SPILL16_256;
  reg Tsfl1_22_V_0;
  integer Tse0SPILL18_256;
  reg Tsfl1_22_V_1;
  reg [63:0] Tsad1_3_V_3;
  reg signed [15:0] Tsad1_3_V_0;
  reg [63:0] Tsad1_3_V_4;
  reg signed [15:0] Tsad1_3_V_1;
  integer Tsad1_3_V_6;
  reg [63:0] Tspr3_2_V_0;
  reg [63:0] Tspr3_2_V_1;
  reg Tspr3_2_V_2;
  reg Tspr3_2_V_3;
  reg Tspr3_2_V_4;
  reg [63:0] Tsa1_SPILL_256;
  reg [63:0] Tssh8_5_V_0;
  reg [63:0] fastspilldup60;
  reg [63:0] Tss8_SPILL_259;
  reg [63:0] Tss8_SPILL_256;
  reg signed [63:0] Tss8_SPILL_258;
  reg [63:0] Tss8_SPILL_257;
  reg signed [15:0] Tsad1_3_V_2;
  reg [63:0] Tspr12_2_V_0;
  reg [63:0] Tspr12_2_V_1;
  reg Tspr12_2_V_2;
  reg Tspr12_2_V_3;
  reg Tspr12_2_V_4;
  reg [63:0] Tssh17_6_V_0;
  reg [63:0] fastspilldup62;
  reg [63:0] Tss17_SPILL_259;
  reg [63:0] Tss17_SPILL_256;
  reg signed [63:0] Tss17_SPILL_258;
  reg [63:0] Tss17_SPILL_257;
  reg [63:0] Tsad1_3_V_5;
  reg [63:0] Tspr21_3_V_0;
  reg [63:0] Tspr21_3_V_1;
  reg Tspr21_3_V_2;
  reg Tspr21_3_V_3;
  reg Tspr21_3_V_4;
  reg signed [15:0] Tsro28_4_V_0;
  reg [63:0] Tsro28_4_V_1;
  reg signed [15:0] Tsro28_4_V_5;
  reg signed [15:0] Tsro28_4_V_6;
  reg [63:0] fastspilldup66;
  reg [63:0] fastspilldup64;
  reg [63:0] Tsr28_SPILL_260;
  reg [63:0] Tsr28_SPILL_256;
  reg signed [63:0] Tsr28_SPILL_258;
  reg [63:0] Tsr28_SPILL_257;
  reg [63:0] Tsr28_SPILL_259;
  reg [63:0] Tsf1SPILL12_256;
  reg Tssu2_4_V_0;
  reg [63:0] Tssu2_4_V_4;
  reg signed [15:0] Tssu2_4_V_1;
  reg [63:0] Tssu2_4_V_5;
  reg signed [15:0] Tssu2_4_V_2;
  integer Tssu2_4_V_7;
  reg [63:0] Tspr27_2_V_0;
  reg [63:0] Tspr27_2_V_1;
  reg Tspr27_2_V_2;
  reg Tspr27_2_V_3;
  reg Tspr27_2_V_4;
  reg [63:0] Tss2_SPILL_256;
  reg [63:0] Tssh32_5_V_0;
  reg [63:0] fastspilldup70;
  reg [63:0] Tss32_SPILL_259;
  reg [63:0] Tss32_SPILL_256;
  reg signed [63:0] Tss32_SPILL_258;
  reg [63:0] Tss32_SPILL_257;
  reg [63:0] Tspr18_2_V_0;
  reg [63:0] Tspr18_2_V_1;
  reg Tspr18_2_V_2;
  reg Tspr18_2_V_3;
  reg Tspr18_2_V_4;
  reg [63:0] Tssh23_6_V_0;
  reg [63:0] fastspilldup68;
  reg [63:0] Tss23_SPILL_259;
  reg [63:0] Tss23_SPILL_256;
  reg signed [63:0] Tss23_SPILL_258;
  reg [63:0] Tss23_SPILL_257;
  reg [63:0] Tspr7_3_V_0;
  reg [63:0] Tspr7_3_V_1;
  reg Tspr7_3_V_2;
  reg Tspr7_3_V_3;
  reg Tspr7_3_V_4;
  reg [63:0] Tssu2_4_V_6;
  reg signed [15:0] Tssu2_4_V_3;
  integer Tsno34_9_V_0;
  reg signed [15:0] Tsro0_16_V_0;
  reg [63:0] Tsro0_16_V_1;
  reg signed [15:0] Tsro0_16_V_5;
  reg signed [15:0] Tsro0_16_V_6;
  reg [63:0] fastspilldup74;
  reg [63:0] fastspilldup72;
  reg [63:0] Tsr0_SPILL_260;
  reg [63:0] Tsr0_SPILL_256;
  reg signed [63:0] Tsr0_SPILL_258;
  reg [63:0] Tsr0_SPILL_257;
  reg [63:0] Tsr0_SPILL_259;
  integer Tsf0SPILL14_256;
  reg Tsfl0_3_V_0;
  reg Tsfl0_3_V_1;
  integer Tsf0SPILL14_257;
  integer Tsf0SPILL14_258;
  reg [63:0] Tdbm0_3_V_2;
  integer fastspilldup76;
  integer Tdb0_SPILL_259;
  integer Tdb0_SPILL_256;
  integer Tdb0_SPILL_258;
  reg [63:0] Tses25_5_V_1;
  reg [63:0] Tsad6_15_V_0;
  reg [63:0] fastspilldup42;
  reg [63:0] Tsa6_SPILL_262;
  reg [63:0] Tsa6_SPILL_257;
  reg signed [63:0] Tsa6_SPILL_260;
  reg [63:0] Tsa6_SPILL_259;
  reg [7:0] A_8_US_CC_SCALbx14_ARA0[258:0];
  reg [63:0] A_64_US_CC_SCALbx12_ARB0[35:0];
  reg [63:0] A_64_US_CC_SCALbx10_ARA0[35:0];
  reg [9:0] xpc10;
 always   @(posedge clk )  begin 
      //Start structure HPR dfsin
      if (reset)  begin 
               Tsfl0_9_V_0 <= 32'd0;
               Tsfl0_9_V_1 <= 32'd0;
               Tsfl0_9_V_2 <= 32'd0;
               Tdsi3_5_V_3 <= 64'd0;
               Tsfl1_7_V_0 <= 32'd0;
               Tsfl1_7_V_1 <= 32'd0;
               Tsfl1_7_V_2 <= 32'd0;
               Tspr4_3_V_2 <= 32'd0;
               Tspr4_3_V_4 <= 32'd0;
               Tspr4_3_V_1 <= 64'd0;
               Tsfl1_18_V_0 <= 32'd0;
               Tsfl1_18_V_1 <= 32'd0;
               Tsfl1_18_V_2 <= 32'd0;
               Tspr2_2_V_2 <= 32'd0;
               Tspr2_2_V_4 <= 32'd0;
               Tspr2_2_V_1 <= 64'd0;
               Tsad1_3_V_0 <= 32'd0;
               Tsad1_3_V_1 <= 32'd0;
               Tsad1_3_V_6 <= 32'd0;
               Tspr3_2_V_2 <= 32'd0;
               Tspr3_2_V_4 <= 32'd0;
               Tspr3_2_V_1 <= 64'd0;
               Tsfl0_3_V_0 <= 32'd0;
               Tdb0_SPILL_259 <= 32'd0;
               fastspilldup76 <= 32'd0;
               Tdb0_SPILL_258 <= 32'd0;
               Tdb0_SPILL_256 <= 32'd0;
               Tdbm0_3_V_1 <= 32'd0;
               done <= 32'd0;
               Tdbm0_3_V_0 <= 32'd0;
               Tsfl0_3_V_1 <= 32'd0;
               Tsf0SPILL14_257 <= 32'd0;
               Tsf0SPILL14_258 <= 32'd0;
               Tsf0SPILL14_256 <= 32'd0;
               Tdbm0_3_V_2 <= 64'd0;
               dfsin_gloops <= 32'd0;
               Tspr3_2_V_0 <= 64'd0;
               Tspr3_2_V_3 <= 32'd0;
               Tsad1_3_V_5 <= 64'd0;
               fastspilldup66 <= 64'd0;
               fastspilldup64 <= 64'd0;
               Tsr28_SPILL_256 <= 64'd0;
               Tsr28_SPILL_260 <= 64'd0;
               Tsr28_SPILL_257 <= 64'd0;
               Tsr28_SPILL_258 <= 64'd0;
               Tsr28_SPILL_259 <= 64'd0;
               Tss8_SPILL_256 <= 64'd0;
               Tss8_SPILL_259 <= 64'd0;
               Tss8_SPILL_257 <= 64'd0;
               Tss8_SPILL_258 <= 64'd0;
               Tsad1_3_V_4 <= 64'd0;
               fastspilldup60 <= 64'd0;
               Tssh8_5_V_0 <= 64'd0;
               Tspr12_2_V_2 <= 32'd0;
               Tspr12_2_V_4 <= 32'd0;
               Tspr12_2_V_1 <= 64'd0;
               Tspr12_2_V_0 <= 64'd0;
               Tspr12_2_V_3 <= 32'd0;
               Tss17_SPILL_256 <= 64'd0;
               Tss17_SPILL_259 <= 64'd0;
               Tss17_SPILL_257 <= 64'd0;
               Tss17_SPILL_258 <= 64'd0;
               fastspilldup62 <= 64'd0;
               Tssh17_6_V_0 <= 64'd0;
               Tspr21_3_V_2 <= 32'd0;
               Tspr21_3_V_4 <= 32'd0;
               Tspr21_3_V_1 <= 64'd0;
               Tsa1_SPILL_256 <= 64'd0;
               Tspr21_3_V_0 <= 64'd0;
               Tspr21_3_V_3 <= 32'd0;
               Tsro28_4_V_0 <= 32'd0;
               Tsad1_3_V_2 <= 32'd0;
               Tsro28_4_V_1 <= 64'd0;
               Tsro28_4_V_5 <= 32'd0;
               Tsro28_4_V_6 <= 32'd0;
               Tssu2_4_V_7 <= 32'd0;
               Tssu2_4_V_2 <= 32'd0;
               Tssu2_4_V_1 <= 32'd0;
               Tspr27_2_V_2 <= 32'd0;
               Tspr27_2_V_4 <= 32'd0;
               Tspr27_2_V_1 <= 64'd0;
               Tspr27_2_V_0 <= 64'd0;
               Tspr27_2_V_3 <= 32'd0;
               Tdsi3_5_V_2 <= 32'd0;
               Tsno34_9_V_0 <= 32'd0;
               Tsro0_16_V_5 <= 32'd0;
               fastspilldup74 <= 64'd0;
               fastspilldup72 <= 64'd0;
               Tsr0_SPILL_256 <= 64'd0;
               Tsr0_SPILL_260 <= 64'd0;
               Tsr0_SPILL_257 <= 64'd0;
               Tsr0_SPILL_258 <= 64'd0;
               Tsr0_SPILL_259 <= 64'd0;
               Tsro0_16_V_6 <= 32'd0;
               Tsro0_16_V_0 <= 32'd0;
               Tsro0_16_V_1 <= 64'd0;
               Tss32_SPILL_256 <= 64'd0;
               Tss32_SPILL_259 <= 64'd0;
               Tss32_SPILL_257 <= 64'd0;
               Tss32_SPILL_258 <= 64'd0;
               fastspilldup70 <= 64'd0;
               Tssh32_5_V_0 <= 64'd0;
               Tspr18_2_V_2 <= 32'd0;
               Tspr18_2_V_4 <= 32'd0;
               Tspr18_2_V_1 <= 64'd0;
               Tspr18_2_V_0 <= 64'd0;
               Tspr18_2_V_3 <= 32'd0;
               Tssu2_4_V_3 <= 32'd0;
               Tss23_SPILL_256 <= 64'd0;
               Tss23_SPILL_259 <= 64'd0;
               Tss23_SPILL_257 <= 64'd0;
               Tss23_SPILL_258 <= 64'd0;
               Tssu2_4_V_5 <= 64'd0;
               fastspilldup68 <= 64'd0;
               Tssh23_6_V_0 <= 64'd0;
               Tspr7_3_V_2 <= 32'd0;
               Tspr7_3_V_4 <= 32'd0;
               Tspr7_3_V_1 <= 64'd0;
               Tspr7_3_V_0 <= 64'd0;
               Tspr7_3_V_3 <= 32'd0;
               Tssu2_4_V_6 <= 64'd0;
               Tss2_SPILL_256 <= 64'd0;
               Tdsi3_5_V_0 <= 64'd0;
               Tsf1SPILL12_256 <= 64'd0;
               Tspr2_2_V_0 <= 64'd0;
               Tspr2_2_V_3 <= 32'd0;
               Tspr5_2_V_2 <= 32'd0;
               Tspr5_2_V_4 <= 32'd0;
               Tspr5_2_V_1 <= 64'd0;
               Tspr5_2_V_0 <= 64'd0;
               Tspr5_2_V_3 <= 32'd0;
               Tsfl1_22_V_0 <= 32'd0;
               Tsfl1_22_V_1 <= 32'd0;
               Tse0SPILL18_256 <= 32'd0;
               Tsad1_3_V_3 <= 64'd0;
               Tssu2_4_V_4 <= 64'd0;
               Tssu2_4_V_0 <= 32'd0;
               Tspr10_2_V_2 <= 32'd0;
               Tspr10_2_V_4 <= 32'd0;
               Tspr10_2_V_1 <= 64'd0;
               Tspr10_2_V_0 <= 64'd0;
               Tspr10_2_V_3 <= 32'd0;
               Tsno18_4_V_0 <= 32'd0;
               Tsfl1_18_V_4 <= 32'd0;
               Tse0SPILL16_256 <= 32'd0;
               Tsno22_4_V_0 <= 32'd0;
               Tsfl1_18_V_3 <= 32'd0;
               Tsfl1_18_V_7 <= 64'd0;
               Tsfl1_18_V_5 <= 32'd0;
               Tses25_5_V_0 <= 64'd0;
               Tsmu26_4_V_1 <= 32'd0;
               Tsmu26_4_V_0 <= 32'd0;
               Tsmu26_4_V_3 <= 32'd0;
               Tsmu26_4_V_2 <= 32'd0;
               Tsmu26_4_V_6 <= 64'd0;
               Tsm26_SPILL_264 <= 64'd0;
               fastspilldup46 <= 64'd0;
               Tsm26_SPILL_259 <= 64'd0;
               Tsm26_SPILL_257 <= 64'd0;
               Tsmu26_4_V_5 <= 64'd0;
               Tsmu26_4_V_7 <= 64'd0;
               Tsm26_SPILL_263 <= 64'd0;
               fastspilldup48 <= 64'd0;
               Tsm26_SPILL_262 <= 64'd0;
               Tsm26_SPILL_260 <= 64'd0;
               Tsfl1_18_V_11 <= 64'd0;
               Tsfl1_18_V_12 <= 64'd0;
               fastspilldup50 <= 64'd0;
               Tss26_SPILL_257 <= 64'd0;
               Tss26_SPILL_262 <= 64'd0;
               Tss26_SPILL_259 <= 64'd0;
               Tss26_SPILL_260 <= 64'd0;
               Tsf1SPILL10_259 <= 64'd0;
               Tsf1SPILL10_257 <= 64'd0;
               Tsro33_4_V_5 <= 32'd0;
               fastspilldup58 <= 64'd0;
               fastspilldup56 <= 64'd0;
               Tsr33_SPILL_256 <= 64'd0;
               Tsr33_SPILL_260 <= 64'd0;
               Tsr33_SPILL_257 <= 64'd0;
               Tsr33_SPILL_258 <= 64'd0;
               Tdsi3_5_V_1 <= 64'd0;
               Tsf1SPILL10_256 <= 64'd0;
               Tsr33_SPILL_259 <= 64'd0;
               Tsro33_4_V_6 <= 32'd0;
               Tsro33_4_V_0 <= 32'd0;
               Tsro33_4_V_1 <= 64'd0;
               Tsad27_13_V_0 <= 64'd0;
               fastspilldup52 <= 64'd0;
               Tsfl1_18_V_10 <= 64'd0;
               Tsa27_SPILL_257 <= 64'd0;
               Tsa27_SPILL_262 <= 64'd0;
               Tsa27_SPILL_259 <= 64'd0;
               Tsa27_SPILL_260 <= 64'd0;
               Tsf1SPILL10_260 <= 64'd0;
               fastspilldup54 <= 64'd0;
               Tsfl1_18_V_9 <= 64'd0;
               Tsmu26_4_V_4 <= 64'd0;
               Tse25_SPILL_257 <= 64'd0;
               Tsmu5_7_V_0 <= 32'd0;
               Tsmu5_7_V_3 <= 32'd0;
               Tsmu5_7_V_2 <= 32'd0;
               Tsmu5_7_V_6 <= 64'd0;
               Tsm5_SPILL_264 <= 64'd0;
               fastspilldup36 <= 64'd0;
               Tsm5_SPILL_259 <= 64'd0;
               Tsm5_SPILL_257 <= 64'd0;
               Tsmu5_7_V_5 <= 64'd0;
               Tsmu5_7_V_7 <= 64'd0;
               Tsm5_SPILL_263 <= 64'd0;
               fastspilldup38 <= 64'd0;
               Tsm5_SPILL_262 <= 64'd0;
               Tsm5_SPILL_260 <= 64'd0;
               Tses25_5_V_4 <= 64'd0;
               Tses25_5_V_5 <= 64'd0;
               fastspilldup40 <= 64'd0;
               Tss5_SPILL_257 <= 64'd0;
               Tss5_SPILL_262 <= 64'd0;
               Tss5_SPILL_259 <= 64'd0;
               Tss5_SPILL_260 <= 64'd0;
               Tse25_SPILL_261 <= 64'd0;
               fastspilldup44 <= 64'd0;
               Tse25_SPILL_260 <= 64'd0;
               Tse25_SPILL_258 <= 64'd0;
               Tsfl1_18_V_8 <= 64'd0;
               Tses25_5_V_1 <= 64'd0;
               Tsad6_15_V_0 <= 64'd0;
               fastspilldup42 <= 64'd0;
               Tses25_5_V_3 <= 64'd0;
               Tsa6_SPILL_257 <= 64'd0;
               Tsa6_SPILL_262 <= 64'd0;
               Tsa6_SPILL_259 <= 64'd0;
               Tsa6_SPILL_260 <= 64'd0;
               Tses25_5_V_2 <= 64'd0;
               Tsmu5_7_V_4 <= 64'd0;
               Tsmu5_7_V_1 <= 32'd0;
               Tses25_5_V_6 <= 64'd0;
               Tsi1_SPILL_257 <= 32'd0;
               Tsco5_4_V_1 <= 32'd0;
               Tsin1_17_V_3 <= 32'd0;
               Tsp5_SPILL_256 <= 64'd0;
               Tsin1_17_V_2 <= 64'd0;
               Tsco5_4_V_0 <= 32'd0;
               Tsin1_17_V_1 <= 32'd0;
               Tsfl1_7_V_3 <= 32'd0;
               Tsfl1_18_V_6 <= 64'd0;
               Tsfl1_7_V_4 <= 32'd0;
               Tsfl1_7_V_6 <= 64'd0;
               Tsfl1_7_V_7 <= 64'd0;
               fastspilldup26 <= 64'd0;
               fastspilldup28 <= 64'd0;
               Tsfl1_7_V_9 <= 64'd0;
               Tsf1_SPILL_260 <= 64'd0;
               fastspilldup30 <= 64'd0;
               Tsf1_SPILL_259 <= 64'd0;
               Tsf1_SPILL_257 <= 64'd0;
               Tsfl1_7_V_5 <= 32'd0;
               fastspilldup34 <= 64'd0;
               fastspilldup32 <= 64'd0;
               Tsi1_SPILL_256 <= 64'd0;
               Tsin1_17_V_0 <= 32'd0;
               Tsf1_SPILL_256 <= 64'd0;
               Tsfl1_7_V_8 <= 64'd0;
               Tspr4_3_V_0 <= 64'd0;
               Tspr4_3_V_3 <= 32'd0;
               Tsf0SPILL10_256 <= 32'd0;
               Tspr11_2_V_2 <= 32'd0;
               Tsf0SPILL12_256 <= 32'd0;
               Tspr11_2_V_4 <= 32'd0;
               Tspr11_2_V_1 <= 64'd0;
               Tspr11_2_V_0 <= 64'd0;
               Tspr11_2_V_3 <= 32'd0;
               Tsno19_4_V_0 <= 32'd0;
               Tsfl0_9_V_3 <= 32'd0;
               Tsco0_2_V_0 <= 64'd0;
               Tsco3_7_V_1 <= 32'd0;
               Tsco0_2_V_1 <= 32'd0;
               Tsno23_4_V_0 <= 32'd0;
               Tsfl0_9_V_4 <= 32'd0;
               Tsfl0_9_V_6 <= 64'd0;
               Tsfl0_9_V_7 <= 64'd0;
               Tsmu24_24_V_1 <= 32'd0;
               Tsmu24_24_V_0 <= 32'd0;
               Tsmu24_24_V_3 <= 32'd0;
               Tsmu24_24_V_2 <= 32'd0;
               Tsmu24_24_V_6 <= 64'd0;
               Tsm24_SPILL_264 <= 64'd0;
               fastspilldup16 <= 64'd0;
               Tsm24_SPILL_259 <= 64'd0;
               Tsm24_SPILL_257 <= 64'd0;
               Tsmu24_24_V_5 <= 64'd0;
               Tsmu24_24_V_7 <= 64'd0;
               Tsm24_SPILL_263 <= 64'd0;
               fastspilldup18 <= 64'd0;
               Tsm24_SPILL_262 <= 64'd0;
               Tsm24_SPILL_260 <= 64'd0;
               Tsfl0_9_V_9 <= 64'd0;
               Tsf0_SPILL_260 <= 64'd0;
               fastspilldup20 <= 64'd0;
               Tsf0_SPILL_259 <= 64'd0;
               Tsf0_SPILL_257 <= 64'd0;
               Tsfl0_9_V_5 <= 32'd0;
               Tsro29_4_V_5 <= 32'd0;
               fastspilldup24 <= 64'd0;
               Tss18_SPILL_260 <= 64'd0;
               fastspilldup22 <= 64'd0;
               Tsr29_SPILL_256 <= 64'd0;
               Tsr29_SPILL_260 <= 64'd0;
               Tsr29_SPILL_257 <= 64'd0;
               Tsr29_SPILL_258 <= 64'd0;
               Tsp27_SPILL_256 <= 64'd0;
               Tsfl0_10_V_0 <= 64'd0;
               Tsf0_SPILL_256 <= 64'd0;
               Tsr29_SPILL_259 <= 64'd0;
               Tss18_SPILL_256 <= 64'd0;
               Tss18_SPILL_259 <= 64'd0;
               Tss18_SPILL_257 <= 64'd0;
               Tss18_SPILL_258 <= 64'd0;
               Tsro29_4_V_6 <= 32'd0;
               Tsro29_4_V_0 <= 32'd0;
               Tsro29_4_V_1 <= 64'd0;
               Tssh18_7_V_0 <= 64'd0;
               Tsfl0_9_V_8 <= 64'd0;
               Tsmu24_24_V_4 <= 64'd0;
               xpc10 <= 32'd0;
               Tsco3_7_V_0 <= 32'd0;
               end 
               else  begin 
              
              case (xpc10)
                  10'sd171/*171:xpc10*/: $display("dfsin: Testbench start");

                  10'sd250/*250:xpc10*/: $display("Test: input=%H expected=%H output=%H ", A_64_US_CC_SCALbx12_ARB0[Tdbm0_3_V_1], A_64_US_CC_SCALbx10_ARA0
                  [Tdbm0_3_V_1], Tdbm0_3_V_2);
              endcase
              if ((32'sd0/*0:USA176*/!=(Tdbm0_3_V_2^A_64_US_CC_SCALbx10_ARA0[Tdbm0_3_V_1])) && (xpc10==10'sd251/*251:xpc10*/)) $display("   hamming error=%H"
                  , Tdbm0_3_V_2^A_64_US_CC_SCALbx10_ARA0[Tdbm0_3_V_1]);
                  
              case (xpc10)
                  10'sd253/*253:xpc10*/:  begin 
                      if ((Tdbm0_3_V_0==32'sd36/*36:Tdbm0.3_V_0*/) && (Tdbm0_3_V_1>=32'sd36))  begin 
                              $display("Result: %1d/%1d", Tdbm0_3_V_0, 32'sd36);
                              $display("RESULT: PASS");
                               end 
                              if ((Tdbm0_3_V_0!=32'sd36/*36:Tdbm0.3_V_0*/) && (Tdbm0_3_V_1>=32'sd36))  begin 
                              $display("Result: %1d/%1d", Tdbm0_3_V_0, 32'sd36);
                              $display("RESULT: FAIL");
                               end 
                               end 
                      
                  10'sd254/*254:xpc10*/:  begin 
                      $display("dfsin: Testbench finished");
                      $display("gloops=%1d", dfsin_gloops);
                       end 
                      endcase
              if ((xpc10==10'sd255/*255:xpc10*/)) $finish(32'sd0);
                  if ((xpc10==10'sd256/*256:xpc10*/))  begin 
                      $display("dfsin: Testbench finished");
                      $display("gloops=%1d", dfsin_gloops);
                       end 
                      if (!(!(32'sd2*Tdsi3_5_V_2*(32'sd1+32'sd2*Tdsi3_5_V_2)))) 
                  case (xpc10)
                      10'sd211/*211:xpc10*/:  begin 
                           xpc10 <= 10'sd619/*619:xpc10*/;
                           Tsin1_17_V_0 <= (32'sd2*Tdsi3_5_V_2*(32'sd1+32'sd2*Tdsi3_5_V_2)<32'sd0);
                           end 
                          
                      10'sd633/*633:xpc10*/:  begin 
                           xpc10 <= 10'sd619/*619:xpc10*/;
                           Tsin1_17_V_0 <= (32'sd2*Tdsi3_5_V_2*(32'sd1+32'sd2*Tdsi3_5_V_2)<32'sd0);
                           Tsf1_SPILL_256 <= 64'h_7fff_ffff_ffff_ffff;
                           end 
                          
                      10'sd635/*635:xpc10*/:  begin 
                           xpc10 <= 10'sd619/*619:xpc10*/;
                           Tsin1_17_V_0 <= (32'sd2*Tdsi3_5_V_2*(32'sd1+32'sd2*Tdsi3_5_V_2)<32'sd0);
                           end 
                          
                      10'sd643/*643:xpc10*/:  begin 
                           xpc10 <= 10'sd619/*619:xpc10*/;
                           Tsin1_17_V_0 <= (32'sd2*Tdsi3_5_V_2*(32'sd1+32'sd2*Tdsi3_5_V_2)<32'sd0);
                           end 
                          
                      10'sd646/*646:xpc10*/:  begin 
                           xpc10 <= 10'sd619/*619:xpc10*/;
                           Tsin1_17_V_0 <= (32'sd2*Tdsi3_5_V_2*(32'sd1+32'sd2*Tdsi3_5_V_2)<32'sd0);
                           Tsf1_SPILL_256 <= 64'h_7fff_ffff_ffff_ffff;
                           end 
                          
                      10'sd647/*647:xpc10*/:  begin 
                           xpc10 <= 10'sd619/*619:xpc10*/;
                           Tsin1_17_V_0 <= (32'sd2*Tdsi3_5_V_2*(32'sd1+32'sd2*Tdsi3_5_V_2)<32'sd0);
                           end 
                          
                      10'sd648/*648:xpc10*/:  begin 
                           xpc10 <= 10'sd619/*619:xpc10*/;
                           Tsin1_17_V_0 <= (32'sd2*Tdsi3_5_V_2*(32'sd1+32'sd2*Tdsi3_5_V_2)<32'sd0);
                           end 
                          
                      10'sd659/*659:xpc10*/:  begin 
                           xpc10 <= 10'sd619/*619:xpc10*/;
                           Tsin1_17_V_0 <= (32'sd2*Tdsi3_5_V_2*(32'sd1+32'sd2*Tdsi3_5_V_2)<32'sd0);
                           end 
                          
                      10'sd704/*704:xpc10*/:  begin 
                           xpc10 <= 10'sd619/*619:xpc10*/;
                           Tsin1_17_V_0 <= (32'sd2*Tdsi3_5_V_2*(32'sd1+32'sd2*Tdsi3_5_V_2)<32'sd0);
                           Tsf1_SPILL_256 <= Tsr29_SPILL_259;
                           end 
                          
                      10'sd714/*714:xpc10*/:  begin 
                           xpc10 <= 10'sd619/*619:xpc10*/;
                           Tsin1_17_V_0 <= (32'sd2*Tdsi3_5_V_2*(32'sd1+32'sd2*Tdsi3_5_V_2)<32'sd0);
                           Tsf1_SPILL_256 <= Tsr29_SPILL_259;
                           end 
                          endcase
                   else 
                  case (xpc10)
                      10'sd211/*211:xpc10*/:  begin 
                           xpc10 <= 10'sd212/*212:xpc10*/;
                           Tsfl1_18_V_6 <= 64'shf_ffff_ffff_ffff&Tsf1_SPILL_256;
                           Tsi1_SPILL_256 <= 64'h0;
                           end 
                          
                      10'sd633/*633:xpc10*/:  begin 
                           xpc10 <= 10'sd634/*634:xpc10*/;
                           Tsi1_SPILL_256 <= 64'h0;
                           Tsf1_SPILL_256 <= 64'h_7fff_ffff_ffff_ffff;
                           end 
                          
                      10'sd635/*635:xpc10*/:  begin 
                           xpc10 <= 10'sd212/*212:xpc10*/;
                           Tsfl1_18_V_6 <= 64'shf_ffff_ffff_ffff&Tsf1_SPILL_256;
                           Tsi1_SPILL_256 <= 64'h0;
                           end 
                          
                      10'sd643/*643:xpc10*/:  begin 
                           xpc10 <= 10'sd212/*212:xpc10*/;
                           Tsfl1_18_V_6 <= 64'shf_ffff_ffff_ffff&Tsf1_SPILL_256;
                           Tsi1_SPILL_256 <= 64'h0;
                           end 
                          
                      10'sd646/*646:xpc10*/:  begin 
                           xpc10 <= 10'sd634/*634:xpc10*/;
                           Tsi1_SPILL_256 <= 64'h0;
                           Tsf1_SPILL_256 <= 64'h_7fff_ffff_ffff_ffff;
                           end 
                          
                      10'sd647/*647:xpc10*/:  begin 
                           xpc10 <= 10'sd212/*212:xpc10*/;
                           Tsfl1_18_V_6 <= 64'shf_ffff_ffff_ffff&Tsf1_SPILL_256;
                           Tsi1_SPILL_256 <= 64'h0;
                           end 
                          
                      10'sd648/*648:xpc10*/:  begin 
                           xpc10 <= 10'sd212/*212:xpc10*/;
                           Tsfl1_18_V_6 <= 64'shf_ffff_ffff_ffff&Tsf1_SPILL_256;
                           Tsi1_SPILL_256 <= 64'h0;
                           end 
                          
                      10'sd659/*659:xpc10*/:  begin 
                           xpc10 <= 10'sd212/*212:xpc10*/;
                           Tsfl1_18_V_6 <= 64'shf_ffff_ffff_ffff&Tsf1_SPILL_256;
                           Tsi1_SPILL_256 <= 64'h0;
                           end 
                          
                      10'sd704/*704:xpc10*/:  begin 
                           xpc10 <= 10'sd634/*634:xpc10*/;
                           Tsi1_SPILL_256 <= 64'h0;
                           Tsf1_SPILL_256 <= Tsr29_SPILL_259;
                           end 
                          
                      10'sd714/*714:xpc10*/:  begin 
                           xpc10 <= 10'sd634/*634:xpc10*/;
                           Tsi1_SPILL_256 <= 64'h0;
                           Tsf1_SPILL_256 <= Tsr29_SPILL_259;
                           end 
                          endcase
              if ((64'sh0<(Tdsi3_5_V_0>>32'sd63))) 
                  case (xpc10)
                      10'sd226/*226:xpc10*/:  begin 
                           xpc10 <= 10'sd227/*227:xpc10*/;
                           Tse0SPILL16_256 <= 32'sd1;
                           Tdsi3_5_V_1 <= Tsf1SPILL10_256;
                           end 
                          
                      10'sd460/*460:xpc10*/:  begin 
                           xpc10 <= 10'sd227/*227:xpc10*/;
                           Tse0SPILL16_256 <= 32'sd1;
                           Tdsi3_5_V_1 <= Tsf1SPILL10_256;
                           end 
                          
                      10'sd464/*464:xpc10*/:  begin 
                           xpc10 <= 10'sd465/*465:xpc10*/;
                           Tsfl1_22_V_0 <= 1'h1;
                           Tse0SPILL16_256 <= 32'sd1;
                           end 
                          
                      10'sd467/*467:xpc10*/:  begin 
                           xpc10 <= 10'sd227/*227:xpc10*/;
                           Tse0SPILL16_256 <= 32'sd1;
                           Tdsi3_5_V_1 <= Tsf1SPILL10_256;
                           end 
                          
                      10'sd475/*475:xpc10*/:  begin 
                           xpc10 <= 10'sd227/*227:xpc10*/;
                           Tse0SPILL16_256 <= 32'sd1;
                           Tdsi3_5_V_1 <= Tsf1SPILL10_256;
                           end 
                          
                      10'sd478/*478:xpc10*/:  begin 
                           xpc10 <= 10'sd227/*227:xpc10*/;
                           Tse0SPILL16_256 <= 32'sd1;
                           Tdsi3_5_V_1 <= Tsf1SPILL10_256;
                           end 
                          
                      10'sd481/*481:xpc10*/:  begin 
                           xpc10 <= 10'sd227/*227:xpc10*/;
                           Tse0SPILL16_256 <= 32'sd1;
                           Tdsi3_5_V_1 <= Tsf1SPILL10_256;
                           end 
                          
                      10'sd492/*492:xpc10*/:  begin 
                           xpc10 <= 10'sd227/*227:xpc10*/;
                           Tse0SPILL16_256 <= 32'sd1;
                           Tdsi3_5_V_1 <= Tsf1SPILL10_256;
                           end 
                          endcase
                   else 
                  case (xpc10)
                      10'sd226/*226:xpc10*/:  begin 
                           xpc10 <= 10'sd450/*450:xpc10*/;
                           Tse0SPILL16_256 <= 32'sd0;
                           Tdsi3_5_V_1 <= Tsf1SPILL10_256;
                           end 
                          
                      10'sd460/*460:xpc10*/:  begin 
                           xpc10 <= 10'sd450/*450:xpc10*/;
                           Tse0SPILL16_256 <= 32'sd0;
                           Tdsi3_5_V_1 <= Tsf1SPILL10_256;
                           end 
                          
                      10'sd464/*464:xpc10*/:  begin 
                           xpc10 <= 10'sd465/*465:xpc10*/;
                           Tsfl1_22_V_0 <= 1'h0;
                           Tse0SPILL16_256 <= 32'sd0;
                           end 
                          
                      10'sd467/*467:xpc10*/:  begin 
                           xpc10 <= 10'sd450/*450:xpc10*/;
                           Tse0SPILL16_256 <= 32'sd0;
                           Tdsi3_5_V_1 <= Tsf1SPILL10_256;
                           end 
                          
                      10'sd475/*475:xpc10*/:  begin 
                           xpc10 <= 10'sd450/*450:xpc10*/;
                           Tse0SPILL16_256 <= 32'sd0;
                           Tdsi3_5_V_1 <= Tsf1SPILL10_256;
                           end 
                          
                      10'sd478/*478:xpc10*/:  begin 
                           xpc10 <= 10'sd450/*450:xpc10*/;
                           Tse0SPILL16_256 <= 32'sd0;
                           Tdsi3_5_V_1 <= Tsf1SPILL10_256;
                           end 
                          
                      10'sd481/*481:xpc10*/:  begin 
                           xpc10 <= 10'sd450/*450:xpc10*/;
                           Tse0SPILL16_256 <= 32'sd0;
                           Tdsi3_5_V_1 <= Tsf1SPILL10_256;
                           end 
                          
                      10'sd492/*492:xpc10*/:  begin 
                           xpc10 <= 10'sd450/*450:xpc10*/;
                           Tse0SPILL16_256 <= 32'sd0;
                           Tdsi3_5_V_1 <= Tsf1SPILL10_256;
                           end 
                          endcase

              case (xpc10)
                  10'sd184/*184:xpc10*/:  begin 
                      if ((Tsfl0_9_V_3!=32'sd2047/*2047:Tsfl0.9_V_3*/) && (Tsfl0_9_V_4!=32'sd2047/*2047:Tsfl0.9_V_4*/) && (Tsfl0_9_V_7
                      !=32'sd0/*0:Tsfl0.9_V_7*/) && !Tsfl0_9_V_4 && !(!Tsfl0_9_V_3))  begin 
                               xpc10 <= 10'sd758/*758:xpc10*/;
                               Tsco0_2_V_1 <= 8'h0;
                               Tsco0_2_V_0 <= Tsfl0_9_V_7;
                               end 
                              if ((Tsfl0_9_V_3!=32'sd2047/*2047:Tsfl0.9_V_3*/) && (Tsfl0_9_V_6!=32'sd0/*0:Tsfl0.9_V_6*/) && (Tsfl0_9_V_4
                      !=32'sd2047/*2047:Tsfl0.9_V_4*/) && !Tsfl0_9_V_3)  begin 
                               xpc10 <= 10'sd747/*747:xpc10*/;
                               Tsco0_2_V_1 <= 8'h0;
                               Tsco0_2_V_0 <= Tsfl0_9_V_6;
                               end 
                              if ((Tsfl0_9_V_3!=32'sd2047/*2047:Tsfl0.9_V_3*/) && (Tsfl0_9_V_4!=32'sd2047/*2047:Tsfl0.9_V_4*/) && !(!Tsfl0_9_V_4
                      ) && !(!Tsfl0_9_V_3))  begin 
                               xpc10 <= 10'sd768/*768:xpc10*/;
                               Tsfl0_9_V_5 <= rtl_signed_bitextract0(-16'sd1023+Tsfl0_9_V_3+Tsfl0_9_V_4);
                               end 
                              if ((Tsfl0_9_V_3!=32'sd2047/*2047:Tsfl0.9_V_3*/) && (Tsfl0_9_V_4!=32'sd2047/*2047:Tsfl0.9_V_4*/) && (Tsfl0_9_V_7
                      ==32'sd0/*0:Tsfl0.9_V_7*/) && !Tsfl0_9_V_4 && !Tsfl0_9_V_2 && !(!Tsfl0_9_V_3))  begin 
                               xpc10 <= 10'sd757/*757:xpc10*/;
                               Tsf0_SPILL_256 <= 64'h0;
                               end 
                              if ((Tsfl0_9_V_3!=32'sd2047/*2047:Tsfl0.9_V_3*/) && (Tsfl0_9_V_4!=32'sd2047/*2047:Tsfl0.9_V_4*/) && (Tsfl0_9_V_7
                      ==32'sd0/*0:Tsfl0.9_V_7*/) && !Tsfl0_9_V_4 && Tsfl0_9_V_2 && !(!Tsfl0_9_V_3))  begin 
                               xpc10 <= 10'sd757/*757:xpc10*/;
                               Tsf0_SPILL_256 <= 64'h_8000_0000_0000_0000;
                               end 
                              if ((Tsfl0_9_V_3!=32'sd2047/*2047:Tsfl0.9_V_3*/) && (Tsfl0_9_V_6==32'sd0/*0:Tsfl0.9_V_6*/) && (Tsfl0_9_V_4
                      !=32'sd2047/*2047:Tsfl0.9_V_4*/) && !Tsfl0_9_V_2 && !Tsfl0_9_V_3)  begin 
                               xpc10 <= 10'sd746/*746:xpc10*/;
                               Tsf0_SPILL_256 <= 64'h0;
                               end 
                              if ((Tsfl0_9_V_3!=32'sd2047/*2047:Tsfl0.9_V_3*/) && (Tsfl0_9_V_6==32'sd0/*0:Tsfl0.9_V_6*/) && (Tsfl0_9_V_4
                      !=32'sd2047/*2047:Tsfl0.9_V_4*/) && Tsfl0_9_V_2 && !Tsfl0_9_V_3)  begin 
                               xpc10 <= 10'sd746/*746:xpc10*/;
                               Tsf0_SPILL_256 <= 64'h_8000_0000_0000_0000;
                               end 
                              if ((Tsfl0_9_V_3!=32'sd2047/*2047:Tsfl0.9_V_3*/) && (Tsfl0_9_V_4==32'sd2047/*2047:Tsfl0.9_V_4*/) && (Tsfl0_9_V_7
                      ==32'sd0/*0:Tsfl0.9_V_7*/) && !Tsfl0_9_V_2 && !(!Tsfl0_9_V_3))  begin 
                               xpc10 <= 10'sd745/*745:xpc10*/;
                               Tsf0_SPILL_256 <= 64'h_7ff0_0000_0000_0000;
                               end 
                              if ((Tsfl0_9_V_3!=32'sd2047/*2047:Tsfl0.9_V_3*/) && (Tsfl0_9_V_4==32'sd2047/*2047:Tsfl0.9_V_4*/) && (Tsfl0_9_V_7
                      ==32'sd0/*0:Tsfl0.9_V_7*/) && Tsfl0_9_V_2 && !(!Tsfl0_9_V_3))  begin 
                               xpc10 <= 10'sd745/*745:xpc10*/;
                               Tsf0_SPILL_256 <= 64'h_fff0_0000_0000_0000;
                               end 
                              if ((Tsfl0_9_V_3!=32'sd2047/*2047:Tsfl0.9_V_3*/) && (Tsfl0_9_V_6!=32'sd0/*0:Tsfl0.9_V_6*/) && (Tsfl0_9_V_4
                      ==32'sd2047/*2047:Tsfl0.9_V_4*/) && (Tsfl0_9_V_7==32'sd0/*0:Tsfl0.9_V_7*/) && !Tsfl0_9_V_2 && !Tsfl0_9_V_3)  begin 
                               xpc10 <= 10'sd745/*745:xpc10*/;
                               Tsf0_SPILL_256 <= 64'h_7ff0_0000_0000_0000;
                               end 
                              if ((Tsfl0_9_V_3!=32'sd2047/*2047:Tsfl0.9_V_3*/) && (Tsfl0_9_V_6!=32'sd0/*0:Tsfl0.9_V_6*/) && (Tsfl0_9_V_4
                      ==32'sd2047/*2047:Tsfl0.9_V_4*/) && (Tsfl0_9_V_7==32'sd0/*0:Tsfl0.9_V_7*/) && Tsfl0_9_V_2 && !Tsfl0_9_V_3)  begin 
                               xpc10 <= 10'sd745/*745:xpc10*/;
                               Tsf0_SPILL_256 <= 64'h_fff0_0000_0000_0000;
                               end 
                              if ((Tsfl0_9_V_3!=32'sd2047/*2047:Tsfl0.9_V_3*/) && (Tsfl0_9_V_4==32'sd2047/*2047:Tsfl0.9_V_4*/) && (Tsfl0_9_V_7
                      !=32'sd0/*0:Tsfl0.9_V_7*/))  begin 
                               xpc10 <= 10'sd733/*733:xpc10*/;
                               Tspr11_2_V_0 <= $unsigned(A_64_US_CC_SCALbx12_ARB0[Tdbm0_3_V_1]);
                               end 
                              if ((Tsfl0_9_V_3==32'sd2047/*2047:Tsfl0.9_V_3*/) && (Tsfl0_9_V_6!=32'sd0/*0:Tsfl0.9_V_6*/))  begin 
                               xpc10 <= 10'sd185/*185:xpc10*/;
                               Tspr4_3_V_0 <= $unsigned(A_64_US_CC_SCALbx12_ARB0[Tdbm0_3_V_1]);
                               end 
                              if ((Tsfl0_9_V_3==32'sd2047/*2047:Tsfl0.9_V_3*/) && (Tsfl0_9_V_6==32'sd0/*0:Tsfl0.9_V_6*/) && (Tsfl0_9_V_4
                      !=32'sd2047/*2047:Tsfl0.9_V_4*/) && !(!Tsfl0_9_V_4) && !Tsfl0_9_V_2)  begin 
                               xpc10 <= 10'sd732/*732:xpc10*/;
                               Tsf0_SPILL_256 <= 64'h_7ff0_0000_0000_0000;
                               end 
                              if ((Tsfl0_9_V_3==32'sd2047/*2047:Tsfl0.9_V_3*/) && (Tsfl0_9_V_6==32'sd0/*0:Tsfl0.9_V_6*/) && (Tsfl0_9_V_4
                      !=32'sd2047/*2047:Tsfl0.9_V_4*/) && !(!Tsfl0_9_V_4) && Tsfl0_9_V_2)  begin 
                               xpc10 <= 10'sd732/*732:xpc10*/;
                               Tsf0_SPILL_256 <= 64'h_fff0_0000_0000_0000;
                               end 
                              if ((Tsfl0_9_V_3==32'sd2047/*2047:Tsfl0.9_V_3*/) && (Tsfl0_9_V_6==32'sd0/*0:Tsfl0.9_V_6*/) && (Tsfl0_9_V_4
                      !=32'sd2047/*2047:Tsfl0.9_V_4*/) && (Tsfl0_9_V_7!=32'sd0/*0:Tsfl0.9_V_7*/) && !Tsfl0_9_V_4 && !Tsfl0_9_V_2)  begin 
                               xpc10 <= 10'sd732/*732:xpc10*/;
                               Tsf0_SPILL_256 <= 64'h_7ff0_0000_0000_0000;
                               end 
                              if ((Tsfl0_9_V_3==32'sd2047/*2047:Tsfl0.9_V_3*/) && (Tsfl0_9_V_6==32'sd0/*0:Tsfl0.9_V_6*/) && (Tsfl0_9_V_4
                      !=32'sd2047/*2047:Tsfl0.9_V_4*/) && (Tsfl0_9_V_7!=32'sd0/*0:Tsfl0.9_V_7*/) && !Tsfl0_9_V_4 && Tsfl0_9_V_2)  begin 
                               xpc10 <= 10'sd732/*732:xpc10*/;
                               Tsf0_SPILL_256 <= 64'h_fff0_0000_0000_0000;
                               end 
                              if ((Tsfl0_9_V_3==32'sd2047/*2047:Tsfl0.9_V_3*/) && (Tsfl0_9_V_6==32'sd0/*0:Tsfl0.9_V_6*/) && (Tsfl0_9_V_4
                      ==32'sd2047/*2047:Tsfl0.9_V_4*/) && (Tsfl0_9_V_7==32'sd0/*0:Tsfl0.9_V_7*/) && !(!Tsfl0_9_V_4) && !Tsfl0_9_V_2) 
                       begin 
                               xpc10 <= 10'sd732/*732:xpc10*/;
                               Tsf0_SPILL_256 <= 64'h_7ff0_0000_0000_0000;
                               end 
                              if ((Tsfl0_9_V_3==32'sd2047/*2047:Tsfl0.9_V_3*/) && (Tsfl0_9_V_6==32'sd0/*0:Tsfl0.9_V_6*/) && (Tsfl0_9_V_4
                      ==32'sd2047/*2047:Tsfl0.9_V_4*/) && (Tsfl0_9_V_7==32'sd0/*0:Tsfl0.9_V_7*/) && !(!Tsfl0_9_V_4) && Tsfl0_9_V_2)  begin 
                               xpc10 <= 10'sd732/*732:xpc10*/;
                               Tsf0_SPILL_256 <= 64'h_fff0_0000_0000_0000;
                               end 
                              if ((Tsfl0_9_V_3==32'sd2047/*2047:Tsfl0.9_V_3*/) && (Tsfl0_9_V_6==32'sd0/*0:Tsfl0.9_V_6*/) && (Tsfl0_9_V_4
                      ==32'sd2047/*2047:Tsfl0.9_V_4*/) && (Tsfl0_9_V_7!=32'sd0/*0:Tsfl0.9_V_7*/))  begin 
                               xpc10 <= 10'sd185/*185:xpc10*/;
                               Tspr4_3_V_0 <= $unsigned(A_64_US_CC_SCALbx12_ARB0[Tdbm0_3_V_1]);
                               end 
                              if ((Tsfl0_9_V_3==32'sd2047/*2047:Tsfl0.9_V_3*/) && (Tsfl0_9_V_6==32'sd0/*0:Tsfl0.9_V_6*/) && (Tsfl0_9_V_4
                      ==32'sd2047/*2047:Tsfl0.9_V_4*/) && (Tsfl0_9_V_7==32'sd0/*0:Tsfl0.9_V_7*/) && !Tsfl0_9_V_4)  xpc10 <= 10'sd731/*731:xpc10*/;
                          if ((Tsfl0_9_V_3==32'sd2047/*2047:Tsfl0.9_V_3*/) && (Tsfl0_9_V_6==32'sd0/*0:Tsfl0.9_V_6*/) && (Tsfl0_9_V_4!=
                      32'sd2047/*2047:Tsfl0.9_V_4*/) && (Tsfl0_9_V_7==32'sd0/*0:Tsfl0.9_V_7*/) && !Tsfl0_9_V_4)  xpc10 <= 10'sd731/*731:xpc10*/;
                          if ((Tsfl0_9_V_3!=32'sd2047/*2047:Tsfl0.9_V_3*/) && (Tsfl0_9_V_6==32'sd0/*0:Tsfl0.9_V_6*/) && (Tsfl0_9_V_4==
                      32'sd2047/*2047:Tsfl0.9_V_4*/) && (Tsfl0_9_V_7==32'sd0/*0:Tsfl0.9_V_7*/) && !Tsfl0_9_V_3)  xpc10 <= 10'sd744/*744:xpc10*/;
                           end 
                      
                  10'sd203/*203:xpc10*/:  begin 
                      if ((Tsfl1_7_V_3!=32'sd2047/*2047:Tsfl1.7_V_3*/) && (Tsfl1_7_V_4!=32'sd2047/*2047:Tsfl1.7_V_4*/) && (Tsfl1_7_V_7
                      !=32'sd0/*0:Tsfl1.7_V_7*/) && !Tsfl1_7_V_4 && !(!Tsfl1_7_V_3))  begin 
                               xpc10 <= 10'sd660/*660:xpc10*/;
                               Tsco0_2_V_1 <= 8'h0;
                               Tsco0_2_V_0 <= Tsfl1_7_V_7;
                               end 
                              if ((Tsfl1_7_V_3!=32'sd2047/*2047:Tsfl1.7_V_3*/) && (Tsfl1_7_V_6!=32'sd0/*0:Tsfl1.7_V_6*/) && (Tsfl1_7_V_4
                      !=32'sd2047/*2047:Tsfl1.7_V_4*/) && !Tsfl1_7_V_3)  begin 
                               xpc10 <= 10'sd649/*649:xpc10*/;
                               Tsco0_2_V_1 <= 8'h0;
                               Tsco0_2_V_0 <= Tsfl1_7_V_6;
                               end 
                              if ((Tsfl1_7_V_3!=32'sd2047/*2047:Tsfl1.7_V_3*/) && (Tsfl1_7_V_4==32'sd2047/*2047:Tsfl1.7_V_4*/) && (Tsfl1_7_V_7
                      !=32'sd0/*0:Tsfl1.7_V_7*/))  begin 
                               xpc10 <= 10'sd636/*636:xpc10*/;
                               Tspr11_2_V_1 <= Tdsi3_5_V_3;
                               Tspr11_2_V_0 <= Tdsi3_5_V_1;
                               end 
                              if ((Tsfl1_7_V_3==32'sd2047/*2047:Tsfl1.7_V_3*/) && (Tsfl1_7_V_6!=32'sd0/*0:Tsfl1.7_V_6*/))  begin 
                               xpc10 <= 10'sd204/*204:xpc10*/;
                               Tspr4_3_V_1 <= Tdsi3_5_V_3;
                               Tspr4_3_V_0 <= Tdsi3_5_V_1;
                               end 
                              if ((Tsfl1_7_V_3==32'sd2047/*2047:Tsfl1.7_V_3*/) && (Tsfl1_7_V_6==32'sd0/*0:Tsfl1.7_V_6*/) && (Tsfl1_7_V_4
                      ==32'sd2047/*2047:Tsfl1.7_V_4*/) && (Tsfl1_7_V_7!=32'sd0/*0:Tsfl1.7_V_7*/))  begin 
                               xpc10 <= 10'sd204/*204:xpc10*/;
                               Tspr4_3_V_1 <= Tdsi3_5_V_3;
                               Tspr4_3_V_0 <= Tdsi3_5_V_1;
                               end 
                              if ((Tsfl1_7_V_3!=32'sd2047/*2047:Tsfl1.7_V_3*/) && (Tsfl1_7_V_4!=32'sd2047/*2047:Tsfl1.7_V_4*/) && !(!Tsfl1_7_V_4
                      ) && !(!Tsfl1_7_V_3))  begin 
                               xpc10 <= 10'sd670/*670:xpc10*/;
                               Tsfl1_7_V_5 <= rtl_signed_bitextract0(-16'sd1023+Tsfl1_7_V_3+Tsfl1_7_V_4);
                               end 
                              if ((Tsfl1_7_V_3!=32'sd2047/*2047:Tsfl1.7_V_3*/) && (Tsfl1_7_V_4!=32'sd2047/*2047:Tsfl1.7_V_4*/) && (Tsfl1_7_V_7
                      ==32'sd0/*0:Tsfl1.7_V_7*/) && !Tsfl1_7_V_4 && !Tsfl1_7_V_2 && !(!Tsfl1_7_V_3))  begin 
                               xpc10 <= 10'sd659/*659:xpc10*/;
                               Tsf1_SPILL_256 <= 64'h0;
                               end 
                              if ((Tsfl1_7_V_3!=32'sd2047/*2047:Tsfl1.7_V_3*/) && (Tsfl1_7_V_4!=32'sd2047/*2047:Tsfl1.7_V_4*/) && (Tsfl1_7_V_7
                      ==32'sd0/*0:Tsfl1.7_V_7*/) && !Tsfl1_7_V_4 && Tsfl1_7_V_2 && !(!Tsfl1_7_V_3))  begin 
                               xpc10 <= 10'sd659/*659:xpc10*/;
                               Tsf1_SPILL_256 <= 64'h_8000_0000_0000_0000;
                               end 
                              if ((Tsfl1_7_V_3!=32'sd2047/*2047:Tsfl1.7_V_3*/) && (Tsfl1_7_V_6==32'sd0/*0:Tsfl1.7_V_6*/) && (Tsfl1_7_V_4
                      !=32'sd2047/*2047:Tsfl1.7_V_4*/) && !Tsfl1_7_V_2 && !Tsfl1_7_V_3)  begin 
                               xpc10 <= 10'sd648/*648:xpc10*/;
                               Tsf1_SPILL_256 <= 64'h0;
                               end 
                              if ((Tsfl1_7_V_3!=32'sd2047/*2047:Tsfl1.7_V_3*/) && (Tsfl1_7_V_6==32'sd0/*0:Tsfl1.7_V_6*/) && (Tsfl1_7_V_4
                      !=32'sd2047/*2047:Tsfl1.7_V_4*/) && Tsfl1_7_V_2 && !Tsfl1_7_V_3)  begin 
                               xpc10 <= 10'sd648/*648:xpc10*/;
                               Tsf1_SPILL_256 <= 64'h_8000_0000_0000_0000;
                               end 
                              if ((Tsfl1_7_V_3!=32'sd2047/*2047:Tsfl1.7_V_3*/) && (Tsfl1_7_V_4==32'sd2047/*2047:Tsfl1.7_V_4*/) && (Tsfl1_7_V_7
                      ==32'sd0/*0:Tsfl1.7_V_7*/) && !Tsfl1_7_V_2 && !(!Tsfl1_7_V_3))  begin 
                               xpc10 <= 10'sd647/*647:xpc10*/;
                               Tsf1_SPILL_256 <= 64'h_7ff0_0000_0000_0000;
                               end 
                              if ((Tsfl1_7_V_3!=32'sd2047/*2047:Tsfl1.7_V_3*/) && (Tsfl1_7_V_4==32'sd2047/*2047:Tsfl1.7_V_4*/) && (Tsfl1_7_V_7
                      ==32'sd0/*0:Tsfl1.7_V_7*/) && Tsfl1_7_V_2 && !(!Tsfl1_7_V_3))  begin 
                               xpc10 <= 10'sd647/*647:xpc10*/;
                               Tsf1_SPILL_256 <= 64'h_fff0_0000_0000_0000;
                               end 
                              if ((Tsfl1_7_V_3!=32'sd2047/*2047:Tsfl1.7_V_3*/) && (Tsfl1_7_V_6!=32'sd0/*0:Tsfl1.7_V_6*/) && (Tsfl1_7_V_4
                      ==32'sd2047/*2047:Tsfl1.7_V_4*/) && (Tsfl1_7_V_7==32'sd0/*0:Tsfl1.7_V_7*/) && !Tsfl1_7_V_2 && !Tsfl1_7_V_3)  begin 
                               xpc10 <= 10'sd647/*647:xpc10*/;
                               Tsf1_SPILL_256 <= 64'h_7ff0_0000_0000_0000;
                               end 
                              if ((Tsfl1_7_V_3!=32'sd2047/*2047:Tsfl1.7_V_3*/) && (Tsfl1_7_V_6!=32'sd0/*0:Tsfl1.7_V_6*/) && (Tsfl1_7_V_4
                      ==32'sd2047/*2047:Tsfl1.7_V_4*/) && (Tsfl1_7_V_7==32'sd0/*0:Tsfl1.7_V_7*/) && Tsfl1_7_V_2 && !Tsfl1_7_V_3)  begin 
                               xpc10 <= 10'sd647/*647:xpc10*/;
                               Tsf1_SPILL_256 <= 64'h_fff0_0000_0000_0000;
                               end 
                              if ((Tsfl1_7_V_3==32'sd2047/*2047:Tsfl1.7_V_3*/) && (Tsfl1_7_V_6==32'sd0/*0:Tsfl1.7_V_6*/) && (Tsfl1_7_V_4
                      !=32'sd2047/*2047:Tsfl1.7_V_4*/) && !(!Tsfl1_7_V_4) && !Tsfl1_7_V_2)  begin 
                               xpc10 <= 10'sd635/*635:xpc10*/;
                               Tsf1_SPILL_256 <= 64'h_7ff0_0000_0000_0000;
                               end 
                              if ((Tsfl1_7_V_3==32'sd2047/*2047:Tsfl1.7_V_3*/) && (Tsfl1_7_V_6==32'sd0/*0:Tsfl1.7_V_6*/) && (Tsfl1_7_V_4
                      !=32'sd2047/*2047:Tsfl1.7_V_4*/) && !(!Tsfl1_7_V_4) && Tsfl1_7_V_2)  begin 
                               xpc10 <= 10'sd635/*635:xpc10*/;
                               Tsf1_SPILL_256 <= 64'h_fff0_0000_0000_0000;
                               end 
                              if ((Tsfl1_7_V_3==32'sd2047/*2047:Tsfl1.7_V_3*/) && (Tsfl1_7_V_6==32'sd0/*0:Tsfl1.7_V_6*/) && (Tsfl1_7_V_4
                      !=32'sd2047/*2047:Tsfl1.7_V_4*/) && (Tsfl1_7_V_7!=32'sd0/*0:Tsfl1.7_V_7*/) && !Tsfl1_7_V_4 && !Tsfl1_7_V_2)  begin 
                               xpc10 <= 10'sd635/*635:xpc10*/;
                               Tsf1_SPILL_256 <= 64'h_7ff0_0000_0000_0000;
                               end 
                              if ((Tsfl1_7_V_3==32'sd2047/*2047:Tsfl1.7_V_3*/) && (Tsfl1_7_V_6==32'sd0/*0:Tsfl1.7_V_6*/) && (Tsfl1_7_V_4
                      !=32'sd2047/*2047:Tsfl1.7_V_4*/) && (Tsfl1_7_V_7!=32'sd0/*0:Tsfl1.7_V_7*/) && !Tsfl1_7_V_4 && Tsfl1_7_V_2)  begin 
                               xpc10 <= 10'sd635/*635:xpc10*/;
                               Tsf1_SPILL_256 <= 64'h_fff0_0000_0000_0000;
                               end 
                              if ((Tsfl1_7_V_3==32'sd2047/*2047:Tsfl1.7_V_3*/) && (Tsfl1_7_V_6==32'sd0/*0:Tsfl1.7_V_6*/) && (Tsfl1_7_V_4
                      ==32'sd2047/*2047:Tsfl1.7_V_4*/) && (Tsfl1_7_V_7==32'sd0/*0:Tsfl1.7_V_7*/) && !(!Tsfl1_7_V_4) && !Tsfl1_7_V_2) 
                       begin 
                               xpc10 <= 10'sd635/*635:xpc10*/;
                               Tsf1_SPILL_256 <= 64'h_7ff0_0000_0000_0000;
                               end 
                              if ((Tsfl1_7_V_3==32'sd2047/*2047:Tsfl1.7_V_3*/) && (Tsfl1_7_V_6==32'sd0/*0:Tsfl1.7_V_6*/) && (Tsfl1_7_V_4
                      ==32'sd2047/*2047:Tsfl1.7_V_4*/) && (Tsfl1_7_V_7==32'sd0/*0:Tsfl1.7_V_7*/) && !(!Tsfl1_7_V_4) && Tsfl1_7_V_2)  begin 
                               xpc10 <= 10'sd635/*635:xpc10*/;
                               Tsf1_SPILL_256 <= 64'h_fff0_0000_0000_0000;
                               end 
                              if ((Tsfl1_7_V_3==32'sd2047/*2047:Tsfl1.7_V_3*/) && (Tsfl1_7_V_6==32'sd0/*0:Tsfl1.7_V_6*/) && (Tsfl1_7_V_4
                      ==32'sd2047/*2047:Tsfl1.7_V_4*/) && (Tsfl1_7_V_7==32'sd0/*0:Tsfl1.7_V_7*/) && !Tsfl1_7_V_4)  xpc10 <= 10'sd633/*633:xpc10*/;
                          if ((Tsfl1_7_V_3==32'sd2047/*2047:Tsfl1.7_V_3*/) && (Tsfl1_7_V_6==32'sd0/*0:Tsfl1.7_V_6*/) && (Tsfl1_7_V_4!=
                      32'sd2047/*2047:Tsfl1.7_V_4*/) && (Tsfl1_7_V_7==32'sd0/*0:Tsfl1.7_V_7*/) && !Tsfl1_7_V_4)  xpc10 <= 10'sd633/*633:xpc10*/;
                          if ((Tsfl1_7_V_3!=32'sd2047/*2047:Tsfl1.7_V_3*/) && (Tsfl1_7_V_6==32'sd0/*0:Tsfl1.7_V_6*/) && (Tsfl1_7_V_4==
                      32'sd2047/*2047:Tsfl1.7_V_4*/) && (Tsfl1_7_V_7==32'sd0/*0:Tsfl1.7_V_7*/) && !Tsfl1_7_V_3)  xpc10 <= 10'sd646/*646:xpc10*/;
                           end 
                      
                  10'sd235/*235:xpc10*/:  begin 
                      if ((32'sd0>=Tsad1_3_V_6) && (Tsad1_3_V_0==32'sd2047/*2047:Tsad1.3_V_0*/) && (Tsad1_3_V_3!=32'sd0/*0:Tsad1.3_V_3*/) && 
                      (Tsad1_3_V_6>=32'sd0))  begin 
                               xpc10 <= 10'sd330/*330:xpc10*/;
                               Tspr21_3_V_1 <= Tdsi3_5_V_1;
                               Tspr21_3_V_0 <= Tdsi3_5_V_0;
                               end 
                              if ((32'sd0>=Tsad1_3_V_6) && (Tsad1_3_V_0==32'sd2047/*2047:Tsad1.3_V_0*/) && (Tsad1_3_V_3==32'sd0/*0:Tsad1.3_V_3*/) && 
                      (Tsad1_3_V_4==32'sd0/*0:Tsad1.3_V_4*/) && (Tsad1_3_V_6>=32'sd0))  begin 
                               xpc10 <= 10'sd266/*266:xpc10*/;
                               Tsf1SPILL12_256 <= Tdsi3_5_V_0;
                               Tsa1_SPILL_256 <= Tdsi3_5_V_0;
                               end 
                              if ((32'sd0>=Tsad1_3_V_6) && (Tsad1_3_V_0==32'sd2047/*2047:Tsad1.3_V_0*/) && (Tsad1_3_V_3==32'sd0/*0:Tsad1.3_V_3*/) && 
                      (Tsad1_3_V_4!=32'sd0/*0:Tsad1.3_V_4*/) && (Tsad1_3_V_6>=32'sd0))  begin 
                               xpc10 <= 10'sd330/*330:xpc10*/;
                               Tspr21_3_V_1 <= Tdsi3_5_V_1;
                               Tspr21_3_V_0 <= Tdsi3_5_V_0;
                               end 
                              if ((Tsad1_3_V_4!=32'sd0/*0:Tsad1.3_V_4*/) && (Tsad1_3_V_6<32'sd0) && (Tsad1_3_V_1==32'sd2047/*2047:Tsad1.3_V_1*/)) 
                       begin 
                               xpc10 <= 10'sd309/*309:xpc10*/;
                               Tspr12_2_V_1 <= Tdsi3_5_V_1;
                               Tspr12_2_V_0 <= Tdsi3_5_V_0;
                               end 
                              if ((32'sd0<Tsad1_3_V_6) && (Tsad1_3_V_0==32'sd2047/*2047:Tsad1.3_V_0*/) && (Tsad1_3_V_3==32'sd0/*0:Tsad1.3_V_3*/)) 
                       begin 
                               xpc10 <= 10'sd266/*266:xpc10*/;
                               Tsf1SPILL12_256 <= Tdsi3_5_V_0;
                               Tsa1_SPILL_256 <= Tdsi3_5_V_0;
                               end 
                              if ((32'sd0<Tsad1_3_V_6) && (Tsad1_3_V_0==32'sd2047/*2047:Tsad1.3_V_0*/) && (Tsad1_3_V_3!=32'sd0/*0:Tsad1.3_V_3*/)) 
                       begin 
                               xpc10 <= 10'sd236/*236:xpc10*/;
                               Tspr3_2_V_1 <= Tdsi3_5_V_1;
                               Tspr3_2_V_0 <= Tdsi3_5_V_0;
                               end 
                              if ((32'sd0>=Tsad1_3_V_6) && (Tsad1_3_V_0!=32'sd2047/*2047:Tsad1.3_V_0*/) && (Tsad1_3_V_6>=32'sd0) && !(!Tsad1_3_V_0
                      ))  begin 
                               xpc10 <= 10'sd341/*341:xpc10*/;
                               Tsad1_3_V_5 <= 64'sh_4000_0000_0000_0000+Tsad1_3_V_3+Tsad1_3_V_4;
                               end 
                              if (!Tsfl1_22_V_0 && (32'sd0>=Tsad1_3_V_6) && (Tsad1_3_V_0!=32'sd2047/*2047:Tsad1.3_V_0*/) && (Tsad1_3_V_6
                      >=32'sd0) && !Tsad1_3_V_0)  begin 
                               xpc10 <= 10'sd340/*340:xpc10*/;
                               Tsa1_SPILL_256 <= (Tsad1_3_V_3+Tsad1_3_V_4>>32'sd9);
                               end 
                              if (Tsfl1_22_V_0 && (32'sd0>=Tsad1_3_V_6) && (Tsad1_3_V_0!=32'sd2047/*2047:Tsad1.3_V_0*/) && (Tsad1_3_V_6
                      >=32'sd0) && !Tsad1_3_V_0)  begin 
                               xpc10 <= 10'sd340/*340:xpc10*/;
                               Tsa1_SPILL_256 <= 64'sh_8000_0000_0000_0000+(Tsad1_3_V_3+Tsad1_3_V_4>>32'sd9);
                               end 
                              if ((Tsad1_3_V_6<32'sd0) && (Tsad1_3_V_1!=32'sd2047/*2047:Tsad1.3_V_1*/) && !(!Tsad1_3_V_0))  begin 
                               xpc10 <= 10'sd329/*329:xpc10*/;
                               Tsad1_3_V_3 <= 64'sh_2000_0000_0000_0000|Tsad1_3_V_3;
                               end 
                              if ((Tsad1_3_V_6<32'sd0) && (Tsad1_3_V_1!=32'sd2047/*2047:Tsad1.3_V_1*/) && !Tsad1_3_V_0)  begin 
                               xpc10 <= 10'sd320/*320:xpc10*/;
                               Tsad1_3_V_6 <= 32'sd1+Tsad1_3_V_6;
                               end 
                              if (!Tsfl1_22_V_0 && (Tsad1_3_V_4==32'sd0/*0:Tsad1.3_V_4*/) && (Tsad1_3_V_6<32'sd0) && (Tsad1_3_V_1==32'sd2047
                      /*2047:Tsad1.3_V_1*/))  begin 
                               xpc10 <= 10'sd319/*319:xpc10*/;
                               Tsa1_SPILL_256 <= 64'h_7ff0_0000_0000_0000;
                               end 
                              if (Tsfl1_22_V_0 && (Tsad1_3_V_4==32'sd0/*0:Tsad1.3_V_4*/) && (Tsad1_3_V_6<32'sd0) && (Tsad1_3_V_1==32'sd2047
                      /*2047:Tsad1.3_V_1*/))  begin 
                               xpc10 <= 10'sd319/*319:xpc10*/;
                               Tsa1_SPILL_256 <= 64'h_fff0_0000_0000_0000;
                               end 
                              if ((32'sd0<Tsad1_3_V_6) && (Tsad1_3_V_0!=32'sd2047/*2047:Tsad1.3_V_0*/) && !(!Tsad1_3_V_1))  begin 
                               xpc10 <= 10'sd308/*308:xpc10*/;
                               Tsad1_3_V_4 <= 64'sh_2000_0000_0000_0000|Tsad1_3_V_4;
                               end 
                              if ((32'sd0<Tsad1_3_V_6) && (Tsad1_3_V_0!=32'sd2047/*2047:Tsad1.3_V_0*/) && !Tsad1_3_V_1)  begin 
                               xpc10 <= 10'sd267/*267:xpc10*/;
                               Tsad1_3_V_6 <= -32'sd1+Tsad1_3_V_6;
                               end 
                               end 
                      
                  10'sd352/*352:xpc10*/:  begin 
                      if ((32'sd0>=Tssu2_4_V_7) && (Tssu2_4_V_1!=32'sd2047/*2047:Tssu2.4_V_1*/) && (Tssu2_4_V_7>=32'sd0) && !Tssu2_4_V_1
                      )  begin 
                               xpc10 <= 10'sd447/*447:xpc10*/;
                               Tssu2_4_V_2 <= 16'sh1;
                               Tssu2_4_V_1 <= 16'sh1;
                               end 
                              if ((32'sd0>=Tssu2_4_V_7) && (Tssu2_4_V_1==32'sd2047/*2047:Tssu2.4_V_1*/) && (Tssu2_4_V_4!=32'sd0/*0:Tssu2.4_V_4*/) && 
                      (Tssu2_4_V_7>=32'sd0))  begin 
                               xpc10 <= 10'sd436/*436:xpc10*/;
                               Tspr7_3_V_1 <= Tdsi3_5_V_1;
                               Tspr7_3_V_0 <= Tdsi3_5_V_0;
                               end 
                              if ((32'sd0>=Tssu2_4_V_7) && (Tssu2_4_V_1==32'sd2047/*2047:Tssu2.4_V_1*/) && (Tssu2_4_V_4==32'sd0/*0:Tssu2.4_V_4*/) && 
                      (Tssu2_4_V_5!=32'sd0/*0:Tssu2.4_V_5*/) && (Tssu2_4_V_7>=32'sd0))  begin 
                               xpc10 <= 10'sd436/*436:xpc10*/;
                               Tspr7_3_V_1 <= Tdsi3_5_V_1;
                               Tspr7_3_V_0 <= Tdsi3_5_V_0;
                               end 
                              if ((Tssu2_4_V_5!=32'sd0/*0:Tssu2.4_V_5*/) && (Tssu2_4_V_7<32'sd0) && (Tssu2_4_V_2==32'sd2047/*2047:Tssu2.4_V_2*/)) 
                       begin 
                               xpc10 <= 10'sd413/*413:xpc10*/;
                               Tspr18_2_V_1 <= Tdsi3_5_V_1;
                               Tspr18_2_V_0 <= Tdsi3_5_V_0;
                               end 
                              if ((32'sd0<Tssu2_4_V_7) && (Tssu2_4_V_1==32'sd2047/*2047:Tssu2.4_V_1*/) && (Tssu2_4_V_4==32'sd0/*0:Tssu2.4_V_4*/)) 
                       begin 
                               xpc10 <= 10'sd363/*363:xpc10*/;
                               Tsf1SPILL12_256 <= Tdsi3_5_V_0;
                               Tss2_SPILL_256 <= Tdsi3_5_V_0;
                               end 
                              if ((32'sd0<Tssu2_4_V_7) && (Tssu2_4_V_1==32'sd2047/*2047:Tssu2.4_V_1*/) && (Tssu2_4_V_4!=32'sd0/*0:Tssu2.4_V_4*/)) 
                       begin 
                               xpc10 <= 10'sd353/*353:xpc10*/;
                               Tspr27_2_V_1 <= Tdsi3_5_V_1;
                               Tspr27_2_V_0 <= Tdsi3_5_V_0;
                               end 
                              if ((32'sd0>=Tssu2_4_V_7) && (Tssu2_4_V_1!=32'sd2047/*2047:Tssu2.4_V_1*/) && (Tssu2_4_V_7>=32'sd0) && !(!Tssu2_4_V_1
                      ) && (Tssu2_4_V_5>=Tssu2_4_V_4) && (Tssu2_4_V_4>=Tssu2_4_V_5))  begin 
                               xpc10 <= 10'sd448/*448:xpc10*/;
                               Tss2_SPILL_256 <= 64'h0;
                               end 
                              if ((32'sd0>=Tssu2_4_V_7) && (Tssu2_4_V_1!=32'sd2047/*2047:Tssu2.4_V_1*/) && (Tssu2_4_V_7>=32'sd0) && !(!Tssu2_4_V_1
                      ) && (Tssu2_4_V_5>=Tssu2_4_V_4) && (Tssu2_4_V_4<Tssu2_4_V_5))  begin 
                               xpc10 <= 10'sd427/*427:xpc10*/;
                               Tssu2_4_V_6 <= Tssu2_4_V_5+(0-Tssu2_4_V_4);
                               end 
                              if ((32'sd0>=Tssu2_4_V_7) && (Tssu2_4_V_1!=32'sd2047/*2047:Tssu2.4_V_1*/) && (Tssu2_4_V_7>=32'sd0) && !(!Tssu2_4_V_1
                      ) && (Tssu2_4_V_5<Tssu2_4_V_4))  begin 
                               xpc10 <= 10'sd367/*367:xpc10*/;
                               Tssu2_4_V_6 <= Tssu2_4_V_4+(0-Tssu2_4_V_5);
                               end 
                              if ((Tssu2_4_V_7<32'sd0) && (Tssu2_4_V_2!=32'sd2047/*2047:Tssu2.4_V_2*/) && !(!Tssu2_4_V_1))  begin 
                               xpc10 <= 10'sd435/*435:xpc10*/;
                               Tssu2_4_V_4 <= 64'sh_4000_0000_0000_0000|Tssu2_4_V_4;
                               end 
                              if ((Tssu2_4_V_7<32'sd0) && (Tssu2_4_V_2!=32'sd2047/*2047:Tssu2.4_V_2*/) && !Tssu2_4_V_1)  begin 
                               xpc10 <= 10'sd424/*424:xpc10*/;
                               Tssu2_4_V_7 <= 32'sd1+Tssu2_4_V_7;
                               end 
                              if ((Tssu2_4_V_5==32'sd0/*0:Tssu2.4_V_5*/) && (Tssu2_4_V_7<32'sd0) && (Tssu2_4_V_2==32'sd2047/*2047:Tssu2.4_V_2*/) && 
                      (Tssu2_4_V_0!=32'sd0/*0:Tssu2.4_V_0*/))  begin 
                               xpc10 <= 10'sd423/*423:xpc10*/;
                               Tss2_SPILL_256 <= 64'h_7ff0_0000_0000_0000;
                               end 
                              if ((Tssu2_4_V_5==32'sd0/*0:Tssu2.4_V_5*/) && (Tssu2_4_V_7<32'sd0) && (Tssu2_4_V_2==32'sd2047/*2047:Tssu2.4_V_2*/) && 
                      (Tssu2_4_V_0==32'sd0/*0:Tssu2.4_V_0*/))  begin 
                               xpc10 <= 10'sd423/*423:xpc10*/;
                               Tss2_SPILL_256 <= 64'h_fff0_0000_0000_0000;
                               end 
                              if ((32'sd0<Tssu2_4_V_7) && (Tssu2_4_V_1!=32'sd2047/*2047:Tssu2.4_V_1*/) && !(!Tssu2_4_V_2))  begin 
                               xpc10 <= 10'sd412/*412:xpc10*/;
                               Tssu2_4_V_5 <= 64'sh_4000_0000_0000_0000|Tssu2_4_V_5;
                               end 
                              if ((32'sd0<Tssu2_4_V_7) && (Tssu2_4_V_1!=32'sd2047/*2047:Tssu2.4_V_1*/) && !Tssu2_4_V_2)  begin 
                               xpc10 <= 10'sd364/*364:xpc10*/;
                               Tssu2_4_V_7 <= -32'sd1+Tssu2_4_V_7;
                               end 
                              if ((32'sd0>=Tssu2_4_V_7) && (Tssu2_4_V_1==32'sd2047/*2047:Tssu2.4_V_1*/) && (Tssu2_4_V_4==32'sd0/*0:Tssu2.4_V_4*/) && 
                      (Tssu2_4_V_5==32'sd0/*0:Tssu2.4_V_5*/) && (Tssu2_4_V_7>=32'sd0))  xpc10 <= 10'sd446/*446:xpc10*/;
                           end 
                      endcase
              if ((Tsco0_2_V_0<64'sh1_0000_0000)) 
                  case (xpc10)
                      10'sd369/*369:xpc10*/:  begin 
                           xpc10 <= 10'sd370/*370:xpc10*/;
                           Tsco3_7_V_0 <= rtl_unsigned_bitextract1(64'h_ffff_ffff&Tsco0_2_V_0);
                           Tsco0_2_V_1 <= 8'h20;
                           end 
                          
                      10'sd482/*482:xpc10*/:  begin 
                           xpc10 <= 10'sd483/*483:xpc10*/;
                           Tsco3_7_V_0 <= rtl_unsigned_bitextract1(64'h_ffff_ffff&Tsco0_2_V_0);
                           Tsco0_2_V_1 <= 8'h20;
                           end 
                          
                      10'sd493/*493:xpc10*/:  begin 
                           xpc10 <= 10'sd494/*494:xpc10*/;
                           Tsco3_7_V_0 <= rtl_unsigned_bitextract1(64'h_ffff_ffff&Tsco0_2_V_0);
                           Tsco0_2_V_1 <= 8'h20;
                           end 
                          
                      10'sd649/*649:xpc10*/:  begin 
                           xpc10 <= 10'sd650/*650:xpc10*/;
                           Tsco3_7_V_0 <= rtl_unsigned_bitextract1(64'h_ffff_ffff&Tsco0_2_V_0);
                           Tsco0_2_V_1 <= 8'h20;
                           end 
                          
                      10'sd660/*660:xpc10*/:  begin 
                           xpc10 <= 10'sd661/*661:xpc10*/;
                           Tsco3_7_V_0 <= rtl_unsigned_bitextract1(64'h_ffff_ffff&Tsco0_2_V_0);
                           Tsco0_2_V_1 <= 8'h20;
                           end 
                          
                      10'sd747/*747:xpc10*/:  begin 
                           xpc10 <= 10'sd748/*748:xpc10*/;
                           Tsco3_7_V_0 <= rtl_unsigned_bitextract1(64'h_ffff_ffff&Tsco0_2_V_0);
                           Tsco0_2_V_1 <= 8'h20;
                           end 
                          
                      10'sd758/*758:xpc10*/:  begin 
                           xpc10 <= 10'sd759/*759:xpc10*/;
                           Tsco3_7_V_0 <= rtl_unsigned_bitextract1(64'h_ffff_ffff&Tsco0_2_V_0);
                           Tsco0_2_V_1 <= 8'h20;
                           end 
                          endcase
                   else 
                  case (xpc10)
                      10'sd369/*369:xpc10*/:  begin 
                           xpc10 <= 10'sd405/*405:xpc10*/;
                           Tsco0_2_V_0 <= (Tsco0_2_V_0>>32'sd32);
                           end 
                          
                      10'sd482/*482:xpc10*/:  begin 
                           xpc10 <= 10'sd618/*618:xpc10*/;
                           Tsco0_2_V_0 <= (Tsco0_2_V_0>>32'sd32);
                           end 
                          
                      10'sd493/*493:xpc10*/:  begin 
                           xpc10 <= 10'sd617/*617:xpc10*/;
                           Tsco0_2_V_0 <= (Tsco0_2_V_0>>32'sd32);
                           end 
                          
                      10'sd649/*649:xpc10*/:  begin 
                           xpc10 <= 10'sd728/*728:xpc10*/;
                           Tsco0_2_V_0 <= (Tsco0_2_V_0>>32'sd32);
                           end 
                          
                      10'sd660/*660:xpc10*/:  begin 
                           xpc10 <= 10'sd727/*727:xpc10*/;
                           Tsco0_2_V_0 <= (Tsco0_2_V_0>>32'sd32);
                           end 
                          
                      10'sd747/*747:xpc10*/:  begin 
                           xpc10 <= 10'sd826/*826:xpc10*/;
                           Tsco0_2_V_0 <= (Tsco0_2_V_0>>32'sd32);
                           end 
                          
                      10'sd758/*758:xpc10*/:  begin 
                           xpc10 <= 10'sd825/*825:xpc10*/;
                           Tsco0_2_V_0 <= (Tsco0_2_V_0>>32'sd32);
                           end 
                          endcase
              if ((xpc10==10'sd218/*218:xpc10*/))  begin 
                      if ((Tsfl1_18_V_3!=32'sd2047/*2047:Tsfl1.18_V_3*/) && (Tsfl1_18_V_6!=32'sd0/*0:Tsfl1.18_V_6*/) && (Tsfl1_18_V_4
                      !=32'sd2047/*2047:Tsfl1.18_V_4*/) && !(!Tsfl1_18_V_4) && !Tsfl1_18_V_3)  begin 
                               xpc10 <= 10'sd493/*493:xpc10*/;
                               Tsco0_2_V_1 <= 8'h0;
                               Tsco0_2_V_0 <= Tsfl1_18_V_6;
                               end 
                              if ((Tsfl1_18_V_3!=32'sd2047/*2047:Tsfl1.18_V_3*/) && (Tsfl1_18_V_4!=32'sd2047/*2047:Tsfl1.18_V_4*/) && 
                      (Tsfl1_18_V_7!=32'sd0/*0:Tsfl1.18_V_7*/) && !Tsfl1_18_V_4)  begin 
                               xpc10 <= 10'sd482/*482:xpc10*/;
                               Tsco0_2_V_1 <= 8'h0;
                               Tsco0_2_V_0 <= Tsfl1_18_V_7;
                               end 
                              if ((Tsfl1_18_V_3!=32'sd2047/*2047:Tsfl1.18_V_3*/) && (Tsfl1_18_V_4==32'sd2047/*2047:Tsfl1.18_V_4*/) && 
                      (Tsfl1_18_V_7!=32'sd0/*0:Tsfl1.18_V_7*/))  begin 
                               xpc10 <= 10'sd468/*468:xpc10*/;
                               Tspr10_2_V_1 <= Tsi1_SPILL_256;
                               Tspr10_2_V_0 <= Tsf1_SPILL_256;
                               end 
                              if ((Tsfl1_18_V_3==32'sd2047/*2047:Tsfl1.18_V_3*/) && (Tsfl1_18_V_6==32'sd0/*0:Tsfl1.18_V_6*/) && (Tsfl1_18_V_4
                      ==32'sd2047/*2047:Tsfl1.18_V_4*/) && (Tsfl1_18_V_7!=32'sd0/*0:Tsfl1.18_V_7*/))  begin 
                               xpc10 <= 10'sd453/*453:xpc10*/;
                               Tspr5_2_V_1 <= Tsi1_SPILL_256;
                               Tspr5_2_V_0 <= Tsf1_SPILL_256;
                               end 
                              if ((Tsfl1_18_V_3==32'sd2047/*2047:Tsfl1.18_V_3*/) && (Tsfl1_18_V_6!=32'sd0/*0:Tsfl1.18_V_6*/))  begin 
                               xpc10 <= 10'sd219/*219:xpc10*/;
                               Tspr2_2_V_1 <= Tsi1_SPILL_256;
                               Tspr2_2_V_0 <= Tsf1_SPILL_256;
                               end 
                              if ((Tsfl1_18_V_3!=32'sd2047/*2047:Tsfl1.18_V_3*/) && (Tsfl1_18_V_4!=32'sd2047/*2047:Tsfl1.18_V_4*/) && 
                      !(!Tsfl1_18_V_4) && !(!Tsfl1_18_V_3))  begin 
                               xpc10 <= 10'sd503/*503:xpc10*/;
                               Tsfl1_18_V_5 <= rtl_signed_bitextract0(rtl_sign_extend2(16'sd1021)+rtl_sign_extend2(Tsfl1_18_V_3)+(0-Tsfl1_18_V_4
                              ));

                               end 
                              if ((Tsfl1_18_V_3!=32'sd2047/*2047:Tsfl1.18_V_3*/) && (Tsfl1_18_V_6==32'sd0/*0:Tsfl1.18_V_6*/) && (Tsfl1_18_V_4
                      !=32'sd2047/*2047:Tsfl1.18_V_4*/) && !Tsfl1_18_V_2 && !(!Tsfl1_18_V_4) && !Tsfl1_18_V_3)  begin 
                               xpc10 <= 10'sd492/*492:xpc10*/;
                               Tsf1SPILL10_256 <= 64'h0;
                               end 
                              if ((Tsfl1_18_V_3!=32'sd2047/*2047:Tsfl1.18_V_3*/) && (Tsfl1_18_V_6==32'sd0/*0:Tsfl1.18_V_6*/) && (Tsfl1_18_V_4
                      !=32'sd2047/*2047:Tsfl1.18_V_4*/) && Tsfl1_18_V_2 && !(!Tsfl1_18_V_4) && !Tsfl1_18_V_3)  begin 
                               xpc10 <= 10'sd492/*492:xpc10*/;
                               Tsf1SPILL10_256 <= 64'h_8000_0000_0000_0000;
                               end 
                              if ((Tsfl1_18_V_3!=32'sd2047/*2047:Tsfl1.18_V_3*/) && (Tsfl1_18_V_4==32'sd2047/*2047:Tsfl1.18_V_4*/) && 
                      (Tsfl1_18_V_7==32'sd0/*0:Tsfl1.18_V_7*/) && !Tsfl1_18_V_2)  begin 
                               xpc10 <= 10'sd478/*478:xpc10*/;
                               Tsf1SPILL10_256 <= 64'h0;
                               end 
                              if ((Tsfl1_18_V_3!=32'sd2047/*2047:Tsfl1.18_V_3*/) && (Tsfl1_18_V_4==32'sd2047/*2047:Tsfl1.18_V_4*/) && 
                      (Tsfl1_18_V_7==32'sd0/*0:Tsfl1.18_V_7*/) && Tsfl1_18_V_2)  begin 
                               xpc10 <= 10'sd478/*478:xpc10*/;
                               Tsf1SPILL10_256 <= 64'h_8000_0000_0000_0000;
                               end 
                              if ((Tsfl1_18_V_3==32'sd2047/*2047:Tsfl1.18_V_3*/) && (Tsfl1_18_V_6==32'sd0/*0:Tsfl1.18_V_6*/) && (Tsfl1_18_V_4
                      !=32'sd2047/*2047:Tsfl1.18_V_4*/) && !Tsfl1_18_V_2)  begin 
                               xpc10 <= 10'sd467/*467:xpc10*/;
                               Tsf1SPILL10_256 <= 64'h_7ff0_0000_0000_0000;
                               end 
                              if ((Tsfl1_18_V_3==32'sd2047/*2047:Tsfl1.18_V_3*/) && (Tsfl1_18_V_6==32'sd0/*0:Tsfl1.18_V_6*/) && (Tsfl1_18_V_4
                      !=32'sd2047/*2047:Tsfl1.18_V_4*/) && Tsfl1_18_V_2)  begin 
                               xpc10 <= 10'sd467/*467:xpc10*/;
                               Tsf1SPILL10_256 <= 64'h_fff0_0000_0000_0000;
                               end 
                              if ((Tsfl1_18_V_3==32'sd2047/*2047:Tsfl1.18_V_3*/) && (Tsfl1_18_V_6==32'sd0/*0:Tsfl1.18_V_6*/) && (Tsfl1_18_V_4
                      ==32'sd2047/*2047:Tsfl1.18_V_4*/) && (Tsfl1_18_V_7==32'sd0/*0:Tsfl1.18_V_7*/))  xpc10 <= 10'sd463/*463:xpc10*/;
                          if ((Tsfl1_18_V_3!=32'sd2047/*2047:Tsfl1.18_V_3*/) && (Tsfl1_18_V_6==32'sd0/*0:Tsfl1.18_V_6*/) && (Tsfl1_18_V_4
                      !=32'sd2047/*2047:Tsfl1.18_V_4*/) && (Tsfl1_18_V_7==32'sd0/*0:Tsfl1.18_V_7*/) && !Tsfl1_18_V_4 && !Tsfl1_18_V_3
                      )  xpc10 <= 10'sd479/*479:xpc10*/;
                          if ((!(!Tsfl1_18_V_3)? 1'd1: (Tsfl1_18_V_6!=32'sd0/*0:Tsfl1.18_V_6*/)) && !Tsfl1_18_V_4 && (Tsfl1_18_V_7==32'sd0
                      /*0:Tsfl1.18_V_7*/) && (Tsfl1_18_V_4!=32'sd2047/*2047:Tsfl1.18_V_4*/) && (Tsfl1_18_V_3!=32'sd2047/*2047:Tsfl1.18_V_3*/)) 
                       xpc10 <= 10'sd480/*480:xpc10*/;
                           end 
                      if ((Tsco3_7_V_0<32'sh100_0000)) 
                  case (xpc10)
                      10'sd371/*371:xpc10*/:  begin 
                           xpc10 <= 10'sd372/*372:xpc10*/;
                           Tsco3_7_V_1 <= rtl_unsigned_bitextract3(8'd8+Tsco3_7_V_1);
                           end 
                          
                      10'sd484/*484:xpc10*/:  begin 
                           xpc10 <= 10'sd485/*485:xpc10*/;
                           Tsco3_7_V_1 <= rtl_unsigned_bitextract3(8'd8+Tsco3_7_V_1);
                           end 
                          
                      10'sd495/*495:xpc10*/:  begin 
                           xpc10 <= 10'sd496/*496:xpc10*/;
                           Tsco3_7_V_1 <= rtl_unsigned_bitextract3(8'd8+Tsco3_7_V_1);
                           end 
                          
                      10'sd651/*651:xpc10*/:  begin 
                           xpc10 <= 10'sd652/*652:xpc10*/;
                           Tsco3_7_V_1 <= rtl_unsigned_bitextract3(8'd8+Tsco3_7_V_1);
                           end 
                          
                      10'sd662/*662:xpc10*/:  begin 
                           xpc10 <= 10'sd663/*663:xpc10*/;
                           Tsco3_7_V_1 <= rtl_unsigned_bitextract3(8'd8+Tsco3_7_V_1);
                           end 
                          
                      10'sd749/*749:xpc10*/:  begin 
                           xpc10 <= 10'sd750/*750:xpc10*/;
                           Tsco3_7_V_1 <= rtl_unsigned_bitextract3(8'd8+Tsco3_7_V_1);
                           end 
                          
                      10'sd760/*760:xpc10*/:  begin 
                           xpc10 <= 10'sd761/*761:xpc10*/;
                           Tsco3_7_V_1 <= rtl_unsigned_bitextract3(8'd8+Tsco3_7_V_1);
                           end 
                          endcase
                   else 
                  case (xpc10)
                      10'sd371/*371:xpc10*/:  begin 
                           xpc10 <= 10'sd374/*374:xpc10*/;
                           Tsco3_7_V_1 <= rtl_unsigned_bitextract3(Tsco3_7_V_1+A_8_US_CC_SCALbx14_ARA0[$unsigned((Tsco3_7_V_0>>32'sd24
                          ))]);

                           end 
                          
                      10'sd484/*484:xpc10*/:  begin 
                           xpc10 <= 10'sd487/*487:xpc10*/;
                           Tsco3_7_V_1 <= rtl_unsigned_bitextract3(Tsco3_7_V_1+A_8_US_CC_SCALbx14_ARA0[$unsigned((Tsco3_7_V_0>>32'sd24
                          ))]);

                           end 
                          
                      10'sd495/*495:xpc10*/:  begin 
                           xpc10 <= 10'sd498/*498:xpc10*/;
                           Tsco3_7_V_1 <= rtl_unsigned_bitextract3(Tsco3_7_V_1+A_8_US_CC_SCALbx14_ARA0[$unsigned((Tsco3_7_V_0>>32'sd24
                          ))]);

                           end 
                          
                      10'sd651/*651:xpc10*/:  begin 
                           xpc10 <= 10'sd654/*654:xpc10*/;
                           Tsco3_7_V_1 <= rtl_unsigned_bitextract3(Tsco3_7_V_1+A_8_US_CC_SCALbx14_ARA0[$unsigned((Tsco3_7_V_0>>32'sd24
                          ))]);

                           end 
                          
                      10'sd662/*662:xpc10*/:  begin 
                           xpc10 <= 10'sd665/*665:xpc10*/;
                           Tsco3_7_V_1 <= rtl_unsigned_bitextract3(Tsco3_7_V_1+A_8_US_CC_SCALbx14_ARA0[$unsigned((Tsco3_7_V_0>>32'sd24
                          ))]);

                           end 
                          
                      10'sd749/*749:xpc10*/:  begin 
                           xpc10 <= 10'sd752/*752:xpc10*/;
                           Tsco3_7_V_1 <= rtl_unsigned_bitextract3(Tsco3_7_V_1+A_8_US_CC_SCALbx14_ARA0[$unsigned((Tsco3_7_V_0>>32'sd24
                          ))]);

                           end 
                          
                      10'sd760/*760:xpc10*/:  begin 
                           xpc10 <= 10'sd763/*763:xpc10*/;
                           Tsco3_7_V_1 <= rtl_unsigned_bitextract3(Tsco3_7_V_1+A_8_US_CC_SCALbx14_ARA0[$unsigned((Tsco3_7_V_0>>32'sd24
                          ))]);

                           end 
                          endcase

              case (xpc10)
                  10'sd276/*276:xpc10*/:  begin 
                      if ((Tsro28_4_V_0>=32'sd2045) && (Tsro28_4_V_0<32'sd0))  begin 
                               xpc10 <= 10'sd283/*283:xpc10*/;
                               Tssh18_7_V_0 <= Tsro28_4_V_1;
                               xpc10 <= 10'sd293/*293:xpc10*/;
                               fastspilldup66 <= (Tsro28_4_V_1>>(32'sd63&rtl_signed_bitextract0((0-Tsro28_4_V_0))));
                               xpc10 <= 10'sd298/*298:xpc10*/;
                               Tss18_SPILL_260 <= 64'sh1;
                               xpc10 <= 10'sd300/*300:xpc10*/;
                               Tss18_SPILL_260 <= 64'sh0;
                               end 
                              if ((Tsro28_4_V_0==32'sd2045/*2045:Tsro28.4_V_0*/) && (Tsro28_4_V_0<32'sd0))  begin 
                               xpc10 <= 10'sd283/*283:xpc10*/;
                               Tssh18_7_V_0 <= Tsro28_4_V_1;
                               xpc10 <= 10'sd293/*293:xpc10*/;
                               fastspilldup66 <= (Tsro28_4_V_1>>(32'sd63&rtl_signed_bitextract0((0-Tsro28_4_V_0))));
                               xpc10 <= 10'sd298/*298:xpc10*/;
                               Tss18_SPILL_260 <= 64'sh1;
                               xpc10 <= 10'sd300/*300:xpc10*/;
                               Tss18_SPILL_260 <= 64'sh0;
                               end 
                              if ((32'sd2045>=Tsro28_4_V_0) && (Tsro28_4_V_0==32'sd2045/*2045:Tsro28.4_V_0*/))  begin 
                               xpc10 <= 10'sd277/*277:xpc10*/;
                               xpc10 <= 10'sd287/*287:xpc10*/;
                               xpc10 <= 10'sd288/*288:xpc10*/;
                               Tsro28_4_V_1 <= (Tsro28_4_V_1+rtl_sign_extend4(Tsro28_4_V_5)>>32'sd10);
                               end 
                              if ((Tsro28_4_V_0<32'sd2045) && !Tsro28_4_V_6)  begin 
                               xpc10 <= 10'sd288/*288:xpc10*/;
                               Tsro28_4_V_1 <= (Tsro28_4_V_1+rtl_sign_extend4(Tsro28_4_V_5)>>32'sd10);
                               end 
                              if ((Tsro28_4_V_0>=32'sd2045) && (32'sd2045>=Tsro28_4_V_0) && !Tsro28_4_V_6)  begin 
                               xpc10 <= 10'sd288/*288:xpc10*/;
                               Tsro28_4_V_1 <= (Tsro28_4_V_1+rtl_sign_extend4(Tsro28_4_V_5)>>32'sd10);
                               end 
                              if ((Tsro28_4_V_0>=32'sd2045) && (32'sd2045>=Tsro28_4_V_0) && !(!Tsro28_4_V_6))  xpc10 <= 10'sd287/*287:xpc10*/;
                          if ((Tsro28_4_V_0>=32'sd2045))  xpc10 <= 10'sd277/*277:xpc10*/;
                          if ((Tsro28_4_V_0<32'sd2045) && !(!Tsro28_4_V_6))  xpc10 <= 10'sd287/*287:xpc10*/;
                           end 
                      
                  10'sd380/*380:xpc10*/:  begin 
                      if ((Tsro0_16_V_0>=32'sd2045) && (Tsro0_16_V_0<32'sd0))  begin 
                               xpc10 <= 10'sd387/*387:xpc10*/;
                               Tssh18_7_V_0 <= Tsro0_16_V_1;
                               xpc10 <= 10'sd397/*397:xpc10*/;
                               fastspilldup74 <= (Tsro0_16_V_1>>(32'sd63&rtl_signed_bitextract0((0-Tsro0_16_V_0))));
                               xpc10 <= 10'sd402/*402:xpc10*/;
                               Tss18_SPILL_260 <= 64'sh1;
                               xpc10 <= 10'sd404/*404:xpc10*/;
                               Tss18_SPILL_260 <= 64'sh0;
                               end 
                              if ((Tsro0_16_V_0==32'sd2045/*2045:Tsro0.16_V_0*/) && (Tsro0_16_V_0<32'sd0))  begin 
                               xpc10 <= 10'sd387/*387:xpc10*/;
                               Tssh18_7_V_0 <= Tsro0_16_V_1;
                               xpc10 <= 10'sd397/*397:xpc10*/;
                               fastspilldup74 <= (Tsro0_16_V_1>>(32'sd63&rtl_signed_bitextract0((0-Tsro0_16_V_0))));
                               xpc10 <= 10'sd402/*402:xpc10*/;
                               Tss18_SPILL_260 <= 64'sh1;
                               xpc10 <= 10'sd404/*404:xpc10*/;
                               Tss18_SPILL_260 <= 64'sh0;
                               end 
                              if ((32'sd2045>=Tsro0_16_V_0) && (Tsro0_16_V_0==32'sd2045/*2045:Tsro0.16_V_0*/))  begin 
                               xpc10 <= 10'sd381/*381:xpc10*/;
                               xpc10 <= 10'sd391/*391:xpc10*/;
                               xpc10 <= 10'sd392/*392:xpc10*/;
                               Tsro0_16_V_1 <= (Tsro0_16_V_1+rtl_sign_extend4(Tsro0_16_V_5)>>32'sd10);
                               end 
                              if ((Tsro0_16_V_0<32'sd2045) && !Tsro0_16_V_6)  begin 
                               xpc10 <= 10'sd392/*392:xpc10*/;
                               Tsro0_16_V_1 <= (Tsro0_16_V_1+rtl_sign_extend4(Tsro0_16_V_5)>>32'sd10);
                               end 
                              if ((Tsro0_16_V_0>=32'sd2045) && (32'sd2045>=Tsro0_16_V_0) && !Tsro0_16_V_6)  begin 
                               xpc10 <= 10'sd392/*392:xpc10*/;
                               Tsro0_16_V_1 <= (Tsro0_16_V_1+rtl_sign_extend4(Tsro0_16_V_5)>>32'sd10);
                               end 
                              if ((Tsro0_16_V_0>=32'sd2045) && (32'sd2045>=Tsro0_16_V_0) && !(!Tsro0_16_V_6))  xpc10 <= 10'sd391/*391:xpc10*/;
                          if ((Tsro0_16_V_0>=32'sd2045))  xpc10 <= 10'sd381/*381:xpc10*/;
                          if ((Tsro0_16_V_0<32'sd2045) && !(!Tsro0_16_V_6))  xpc10 <= 10'sd391/*391:xpc10*/;
                           end 
                      
                  10'sd538/*538:xpc10*/:  begin 
                      if ((Tsro33_4_V_0>=32'sd2045) && (Tsro33_4_V_0<32'sd0))  begin 
                               xpc10 <= 10'sd545/*545:xpc10*/;
                               Tssh18_7_V_0 <= Tsro33_4_V_1;
                               xpc10 <= 10'sd555/*555:xpc10*/;
                               fastspilldup58 <= (Tsro33_4_V_1>>(32'sd63&rtl_signed_bitextract0((0-Tsro33_4_V_0))));
                               xpc10 <= 10'sd560/*560:xpc10*/;
                               Tss18_SPILL_260 <= 64'sh1;
                               xpc10 <= 10'sd562/*562:xpc10*/;
                               Tss18_SPILL_260 <= 64'sh0;
                               end 
                              if ((Tsro33_4_V_0==32'sd2045/*2045:Tsro33.4_V_0*/) && (Tsro33_4_V_0<32'sd0))  begin 
                               xpc10 <= 10'sd545/*545:xpc10*/;
                               Tssh18_7_V_0 <= Tsro33_4_V_1;
                               xpc10 <= 10'sd555/*555:xpc10*/;
                               fastspilldup58 <= (Tsro33_4_V_1>>(32'sd63&rtl_signed_bitextract0((0-Tsro33_4_V_0))));
                               xpc10 <= 10'sd560/*560:xpc10*/;
                               Tss18_SPILL_260 <= 64'sh1;
                               xpc10 <= 10'sd562/*562:xpc10*/;
                               Tss18_SPILL_260 <= 64'sh0;
                               end 
                              if ((32'sd2045>=Tsro33_4_V_0) && (Tsro33_4_V_0==32'sd2045/*2045:Tsro33.4_V_0*/))  begin 
                               xpc10 <= 10'sd539/*539:xpc10*/;
                               xpc10 <= 10'sd549/*549:xpc10*/;
                               xpc10 <= 10'sd550/*550:xpc10*/;
                               Tsro33_4_V_1 <= (Tsro33_4_V_1+rtl_sign_extend4(Tsro33_4_V_5)>>32'sd10);
                               end 
                              if ((Tsro33_4_V_0<32'sd2045) && !Tsro33_4_V_6)  begin 
                               xpc10 <= 10'sd550/*550:xpc10*/;
                               Tsro33_4_V_1 <= (Tsro33_4_V_1+rtl_sign_extend4(Tsro33_4_V_5)>>32'sd10);
                               end 
                              if ((Tsro33_4_V_0>=32'sd2045) && (32'sd2045>=Tsro33_4_V_0) && !Tsro33_4_V_6)  begin 
                               xpc10 <= 10'sd550/*550:xpc10*/;
                               Tsro33_4_V_1 <= (Tsro33_4_V_1+rtl_sign_extend4(Tsro33_4_V_5)>>32'sd10);
                               end 
                              if ((Tsro33_4_V_0>=32'sd2045) && (32'sd2045>=Tsro33_4_V_0) && !(!Tsro33_4_V_6))  xpc10 <= 10'sd549/*549:xpc10*/;
                          if ((Tsro33_4_V_0>=32'sd2045))  xpc10 <= 10'sd539/*539:xpc10*/;
                          if ((Tsro33_4_V_0<32'sd2045) && !(!Tsro33_4_V_6))  xpc10 <= 10'sd549/*549:xpc10*/;
                           end 
                      
                  10'sd699/*699:xpc10*/:  begin 
                      if ((Tsro29_4_V_0>=32'sd2045) && (Tsro29_4_V_0<32'sd0))  begin 
                               xpc10 <= 10'sd706/*706:xpc10*/;
                               Tssh18_7_V_0 <= Tsro29_4_V_1;
                               xpc10 <= 10'sd716/*716:xpc10*/;
                               fastspilldup34 <= (Tsro29_4_V_1>>(32'sd63&rtl_signed_bitextract0((0-Tsro29_4_V_0))));
                               xpc10 <= 10'sd721/*721:xpc10*/;
                               Tss18_SPILL_260 <= 64'sh1;
                               xpc10 <= 10'sd723/*723:xpc10*/;
                               Tss18_SPILL_260 <= 64'sh0;
                               end 
                              if ((Tsro29_4_V_0==32'sd2045/*2045:Tsro29.4_V_0*/) && (Tsro29_4_V_0<32'sd0))  begin 
                               xpc10 <= 10'sd706/*706:xpc10*/;
                               Tssh18_7_V_0 <= Tsro29_4_V_1;
                               xpc10 <= 10'sd716/*716:xpc10*/;
                               fastspilldup34 <= (Tsro29_4_V_1>>(32'sd63&rtl_signed_bitextract0((0-Tsro29_4_V_0))));
                               xpc10 <= 10'sd721/*721:xpc10*/;
                               Tss18_SPILL_260 <= 64'sh1;
                               xpc10 <= 10'sd723/*723:xpc10*/;
                               Tss18_SPILL_260 <= 64'sh0;
                               end 
                              if ((32'sd2045>=Tsro29_4_V_0) && (Tsro29_4_V_0==32'sd2045/*2045:Tsro29.4_V_0*/))  begin 
                               xpc10 <= 10'sd700/*700:xpc10*/;
                               xpc10 <= 10'sd710/*710:xpc10*/;
                               xpc10 <= 10'sd711/*711:xpc10*/;
                               Tsro29_4_V_1 <= (Tsro29_4_V_1+rtl_sign_extend4(Tsro29_4_V_5)>>32'sd10);
                               end 
                              if ((Tsro29_4_V_0<32'sd2045) && !Tsro29_4_V_6)  begin 
                               xpc10 <= 10'sd711/*711:xpc10*/;
                               Tsro29_4_V_1 <= (Tsro29_4_V_1+rtl_sign_extend4(Tsro29_4_V_5)>>32'sd10);
                               end 
                              if ((Tsro29_4_V_0>=32'sd2045) && (32'sd2045>=Tsro29_4_V_0) && !Tsro29_4_V_6)  begin 
                               xpc10 <= 10'sd711/*711:xpc10*/;
                               Tsro29_4_V_1 <= (Tsro29_4_V_1+rtl_sign_extend4(Tsro29_4_V_5)>>32'sd10);
                               end 
                              if ((Tsro29_4_V_0<32'sd2045) && !(!Tsro29_4_V_6))  xpc10 <= 10'sd710/*710:xpc10*/;
                          if ((Tsro29_4_V_0>=32'sd2045))  xpc10 <= 10'sd700/*700:xpc10*/;
                          if ((Tsro29_4_V_0>=32'sd2045) && (32'sd2045>=Tsro29_4_V_0) && !(!Tsro29_4_V_6))  xpc10 <= 10'sd710/*710:xpc10*/;
                           end 
                      
                  10'sd797/*797:xpc10*/:  begin 
                      if ((Tsro29_4_V_0>=32'sd2045) && (Tsro29_4_V_0<32'sd0))  begin 
                               xpc10 <= 10'sd804/*804:xpc10*/;
                               Tssh18_7_V_0 <= Tsro29_4_V_1;
                               xpc10 <= 10'sd814/*814:xpc10*/;
                               fastspilldup24 <= (Tsro29_4_V_1>>(32'sd63&rtl_signed_bitextract0((0-Tsro29_4_V_0))));
                               xpc10 <= 10'sd819/*819:xpc10*/;
                               Tss18_SPILL_260 <= 64'sh1;
                               xpc10 <= 10'sd821/*821:xpc10*/;
                               Tss18_SPILL_260 <= 64'sh0;
                               end 
                              if ((Tsro29_4_V_0==32'sd2045/*2045:Tsro29.4_V_0*/) && (Tsro29_4_V_0<32'sd0))  begin 
                               xpc10 <= 10'sd804/*804:xpc10*/;
                               Tssh18_7_V_0 <= Tsro29_4_V_1;
                               xpc10 <= 10'sd814/*814:xpc10*/;
                               fastspilldup24 <= (Tsro29_4_V_1>>(32'sd63&rtl_signed_bitextract0((0-Tsro29_4_V_0))));
                               xpc10 <= 10'sd819/*819:xpc10*/;
                               Tss18_SPILL_260 <= 64'sh1;
                               xpc10 <= 10'sd821/*821:xpc10*/;
                               Tss18_SPILL_260 <= 64'sh0;
                               end 
                              if ((32'sd2045>=Tsro29_4_V_0) && (Tsro29_4_V_0==32'sd2045/*2045:Tsro29.4_V_0*/))  begin 
                               xpc10 <= 10'sd798/*798:xpc10*/;
                               xpc10 <= 10'sd808/*808:xpc10*/;
                               xpc10 <= 10'sd809/*809:xpc10*/;
                               Tsro29_4_V_1 <= (Tsro29_4_V_1+rtl_sign_extend4(Tsro29_4_V_5)>>32'sd10);
                               end 
                              if ((Tsro29_4_V_0<32'sd2045) && !Tsro29_4_V_6)  begin 
                               xpc10 <= 10'sd809/*809:xpc10*/;
                               Tsro29_4_V_1 <= (Tsro29_4_V_1+rtl_sign_extend4(Tsro29_4_V_5)>>32'sd10);
                               end 
                              if ((Tsro29_4_V_0>=32'sd2045) && (32'sd2045>=Tsro29_4_V_0) && !Tsro29_4_V_6)  begin 
                               xpc10 <= 10'sd809/*809:xpc10*/;
                               Tsro29_4_V_1 <= (Tsro29_4_V_1+rtl_sign_extend4(Tsro29_4_V_5)>>32'sd10);
                               end 
                              if ((Tsro29_4_V_0<32'sd2045) && !(!Tsro29_4_V_6))  xpc10 <= 10'sd808/*808:xpc10*/;
                          if ((Tsro29_4_V_0>=32'sd2045))  xpc10 <= 10'sd798/*798:xpc10*/;
                          if ((Tsro29_4_V_0>=32'sd2045) && (32'sd2045>=Tsro29_4_V_0) && !(!Tsro29_4_V_6))  xpc10 <= 10'sd808/*808:xpc10*/;
                           end 
                      endcase
              if ((64'sh0<(Tdsi3_5_V_1>>32'sd63))) 
                  case (xpc10)
                      10'sd198/*198:xpc10*/:  begin 
                           xpc10 <= 10'sd199/*199:xpc10*/;
                           Tsfl1_7_V_0 <= 1'h1;
                           end 
                          
                      10'sd227/*227:xpc10*/:  begin 
                           xpc10 <= 10'sd228/*228:xpc10*/;
                           Tse0SPILL18_256 <= 32'sd1;
                           Tsfl1_22_V_0 <= rtl_unsigned_bitextract5(Tse0SPILL16_256);
                           end 
                          
                      10'sd450/*450:xpc10*/:  begin 
                           xpc10 <= 10'sd228/*228:xpc10*/;
                           Tse0SPILL18_256 <= 32'sd1;
                           Tsfl1_22_V_0 <= rtl_unsigned_bitextract5(Tse0SPILL16_256);
                           end 
                          
                      10'sd465/*465:xpc10*/:  begin 
                           xpc10 <= 10'sd466/*466:xpc10*/;
                           Tsfl1_22_V_1 <= 1'h1;
                           Tse0SPILL18_256 <= 32'sd1;
                           end 
                          endcase
                   else 
                  case (xpc10)
                      10'sd198/*198:xpc10*/:  begin 
                           xpc10 <= 10'sd199/*199:xpc10*/;
                           Tsfl1_7_V_0 <= 1'h0;
                           end 
                          
                      10'sd227/*227:xpc10*/:  begin 
                           xpc10 <= 10'sd449/*449:xpc10*/;
                           Tse0SPILL18_256 <= 32'sd0;
                           Tsfl1_22_V_0 <= rtl_unsigned_bitextract5(Tse0SPILL16_256);
                           end 
                          
                      10'sd450/*450:xpc10*/:  begin 
                           xpc10 <= 10'sd449/*449:xpc10*/;
                           Tse0SPILL18_256 <= 32'sd0;
                           Tsfl1_22_V_0 <= rtl_unsigned_bitextract5(Tse0SPILL16_256);
                           end 
                          
                      10'sd465/*465:xpc10*/:  begin 
                           xpc10 <= 10'sd466/*466:xpc10*/;
                           Tsfl1_22_V_1 <= 1'h0;
                           Tse0SPILL18_256 <= 32'sd0;
                           end 
                          endcase
              if ((Tsco3_7_V_0>=32'sh1_0000) && (Tsco3_7_V_0<32'sh100_0000)) 
                  case (xpc10)
                      10'sd370/*370:xpc10*/:  begin 
                           xpc10 <= 10'sd373/*373:xpc10*/;
                           Tsco3_7_V_0 <= (Tsco3_7_V_0<<32'sd8);
                           Tsco3_7_V_1 <= 8'h8;
                           end 
                          
                      10'sd483/*483:xpc10*/:  begin 
                           xpc10 <= 10'sd486/*486:xpc10*/;
                           Tsco3_7_V_0 <= (Tsco3_7_V_0<<32'sd8);
                           Tsco3_7_V_1 <= 8'h8;
                           end 
                          
                      10'sd494/*494:xpc10*/:  begin 
                           xpc10 <= 10'sd497/*497:xpc10*/;
                           Tsco3_7_V_0 <= (Tsco3_7_V_0<<32'sd8);
                           Tsco3_7_V_1 <= 8'h8;
                           end 
                          
                      10'sd650/*650:xpc10*/:  begin 
                           xpc10 <= 10'sd653/*653:xpc10*/;
                           Tsco3_7_V_0 <= (Tsco3_7_V_0<<32'sd8);
                           Tsco3_7_V_1 <= 8'h8;
                           end 
                          
                      10'sd661/*661:xpc10*/:  begin 
                           xpc10 <= 10'sd664/*664:xpc10*/;
                           Tsco3_7_V_0 <= (Tsco3_7_V_0<<32'sd8);
                           Tsco3_7_V_1 <= 8'h8;
                           end 
                          
                      10'sd748/*748:xpc10*/:  begin 
                           xpc10 <= 10'sd751/*751:xpc10*/;
                           Tsco3_7_V_0 <= (Tsco3_7_V_0<<32'sd8);
                           Tsco3_7_V_1 <= 8'h8;
                           end 
                          
                      10'sd759/*759:xpc10*/:  begin 
                           xpc10 <= 10'sd762/*762:xpc10*/;
                           Tsco3_7_V_0 <= (Tsco3_7_V_0<<32'sd8);
                           Tsco3_7_V_1 <= 8'h8;
                           end 
                          endcase
                  if ((Tsco3_7_V_0<32'sh1_0000)) 
                  case (xpc10)
                      10'sd370/*370:xpc10*/:  begin 
                           xpc10 <= 10'sd371/*371:xpc10*/;
                           Tsco3_7_V_0 <= (Tsco3_7_V_0<<32'sd16);
                           Tsco3_7_V_1 <= 8'h10;
                           end 
                          
                      10'sd483/*483:xpc10*/:  begin 
                           xpc10 <= 10'sd484/*484:xpc10*/;
                           Tsco3_7_V_0 <= (Tsco3_7_V_0<<32'sd16);
                           Tsco3_7_V_1 <= 8'h10;
                           end 
                          
                      10'sd494/*494:xpc10*/:  begin 
                           xpc10 <= 10'sd495/*495:xpc10*/;
                           Tsco3_7_V_0 <= (Tsco3_7_V_0<<32'sd16);
                           Tsco3_7_V_1 <= 8'h10;
                           end 
                          
                      10'sd650/*650:xpc10*/:  begin 
                           xpc10 <= 10'sd651/*651:xpc10*/;
                           Tsco3_7_V_0 <= (Tsco3_7_V_0<<32'sd16);
                           Tsco3_7_V_1 <= 8'h10;
                           end 
                          
                      10'sd661/*661:xpc10*/:  begin 
                           xpc10 <= 10'sd662/*662:xpc10*/;
                           Tsco3_7_V_0 <= (Tsco3_7_V_0<<32'sd16);
                           Tsco3_7_V_1 <= 8'h10;
                           end 
                          
                      10'sd748/*748:xpc10*/:  begin 
                           xpc10 <= 10'sd749/*749:xpc10*/;
                           Tsco3_7_V_0 <= (Tsco3_7_V_0<<32'sd16);
                           Tsco3_7_V_1 <= 8'h10;
                           end 
                          
                      10'sd759/*759:xpc10*/:  begin 
                           xpc10 <= 10'sd760/*760:xpc10*/;
                           Tsco3_7_V_0 <= (Tsco3_7_V_0<<32'sd16);
                           Tsco3_7_V_1 <= 8'h10;
                           end 
                          endcase
                  
              case (xpc10)
                  10'sd392/*392:xpc10*/:  begin 
                      if (!Tssu2_4_V_0 && (Tsro0_16_V_1!=32'sd0/*0:Tsro0.16_V_1*/) && !(32'sd1&(32'sd0/*0:USA164*/==(32'sd512^Tsro0_16_V_6
                      ))))  begin 
                               xpc10 <= 10'sd395/*395:xpc10*/;
                               Tsr0_SPILL_259 <= Tsro0_16_V_1+(rtl_sign_extend4(Tsro0_16_V_0)<<32'sd52);
                               Tsp27_SPILL_256 <= 64'sh0;
                               end 
                              if (Tssu2_4_V_0 && (Tsro0_16_V_1!=32'sd0/*0:Tsro0.16_V_1*/) && !(32'sd1&(32'sd0/*0:USA164*/==(32'sd512^
                      Tsro0_16_V_6))))  begin 
                               xpc10 <= 10'sd395/*395:xpc10*/;
                               Tsr0_SPILL_259 <= 64'sh_8000_0000_0000_0000+Tsro0_16_V_1+(rtl_sign_extend4(Tsro0_16_V_0)<<32'sd52);
                               Tsp27_SPILL_256 <= 64'sh1;
                               end 
                              if (!Tssu2_4_V_0 && (Tsro0_16_V_1==32'sd0/*0:Tsro0.16_V_1*/) && !(32'sd1&(32'sd0/*0:USA164*/==(32'sd512
                      ^Tsro0_16_V_6))))  begin 
                               xpc10 <= 10'sd396/*396:xpc10*/;
                               Tsp27_SPILL_256 <= 64'sh0;
                               Tsro0_16_V_0 <= 16'sh0;
                               end 
                              if (Tssu2_4_V_0 && (Tsro0_16_V_1==32'sd0/*0:Tsro0.16_V_1*/) && !(32'sd1&(32'sd0/*0:USA164*/==(32'sd512^
                      Tsro0_16_V_6))))  begin 
                               xpc10 <= 10'sd394/*394:xpc10*/;
                               Tsp27_SPILL_256 <= 64'sh1;
                               Tsro0_16_V_0 <= 16'sh0;
                               end 
                              if (32'sd1&(32'sd0/*0:USA164*/==(32'sd512^Tsro0_16_V_6)))  begin 
                               xpc10 <= 10'sd393/*393:xpc10*/;
                               Tsro0_16_V_1 <= -64'sh2&Tsro0_16_V_1;
                               end 
                               end 
                      
                  10'sd550/*550:xpc10*/:  begin 
                      if (!Tsfl1_18_V_2 && (Tsro33_4_V_1!=32'sd0/*0:Tsro33.4_V_1*/) && !(32'sd1&(32'sd0/*0:USA76*/==(32'sd512^Tsro33_4_V_6
                      ))))  begin 
                               xpc10 <= 10'sd553/*553:xpc10*/;
                               Tsr33_SPILL_259 <= Tsro33_4_V_1+(rtl_sign_extend4(Tsro33_4_V_0)<<32'sd52);
                               Tsp27_SPILL_256 <= 64'sh0;
                               end 
                              if (Tsfl1_18_V_2 && (Tsro33_4_V_1!=32'sd0/*0:Tsro33.4_V_1*/) && !(32'sd1&(32'sd0/*0:USA76*/==(32'sd512^
                      Tsro33_4_V_6))))  begin 
                               xpc10 <= 10'sd553/*553:xpc10*/;
                               Tsr33_SPILL_259 <= 64'sh_8000_0000_0000_0000+Tsro33_4_V_1+(rtl_sign_extend4(Tsro33_4_V_0)<<32'sd52);
                               Tsp27_SPILL_256 <= 64'sh1;
                               end 
                              if (!Tsfl1_18_V_2 && (Tsro33_4_V_1==32'sd0/*0:Tsro33.4_V_1*/) && !(32'sd1&(32'sd0/*0:USA76*/==(32'sd512
                      ^Tsro33_4_V_6))))  begin 
                               xpc10 <= 10'sd554/*554:xpc10*/;
                               Tsp27_SPILL_256 <= 64'sh0;
                               Tsro33_4_V_0 <= 16'sh0;
                               end 
                              if (Tsfl1_18_V_2 && (Tsro33_4_V_1==32'sd0/*0:Tsro33.4_V_1*/) && !(32'sd1&(32'sd0/*0:USA76*/==(32'sd512^
                      Tsro33_4_V_6))))  begin 
                               xpc10 <= 10'sd552/*552:xpc10*/;
                               Tsp27_SPILL_256 <= 64'sh1;
                               Tsro33_4_V_0 <= 16'sh0;
                               end 
                              if (32'sd1&(32'sd0/*0:USA76*/==(32'sd512^Tsro33_4_V_6)))  begin 
                               xpc10 <= 10'sd551/*551:xpc10*/;
                               Tsro33_4_V_1 <= -64'sh2&Tsro33_4_V_1;
                               end 
                               end 
                      
                  10'sd711/*711:xpc10*/:  begin 
                      if (32'sd1&(32'sd0/*0:USA36*/==(32'sd512^Tsro29_4_V_6)))  begin 
                               xpc10 <= 10'sd712/*712:xpc10*/;
                               Tsro29_4_V_1 <= -64'sh2&Tsro29_4_V_1;
                               end 
                              if ((Tsro29_4_V_1!=32'sd0/*0:Tsro29.4_V_1*/) && !(32'sd1&(32'sd0/*0:USA36*/==(32'sd512^Tsro29_4_V_6))) && 
                      !Tsfl1_7_V_2)  begin 
                               xpc10 <= 10'sd714/*714:xpc10*/;
                               Tsr29_SPILL_259 <= Tsro29_4_V_1+(rtl_sign_extend4(Tsro29_4_V_0)<<32'sd52);
                               Tsp27_SPILL_256 <= 64'sh0;
                               end 
                              if ((Tsro29_4_V_1!=32'sd0/*0:Tsro29.4_V_1*/) && !(32'sd1&(32'sd0/*0:USA36*/==(32'sd512^Tsro29_4_V_6))) && 
                      Tsfl1_7_V_2)  begin 
                               xpc10 <= 10'sd714/*714:xpc10*/;
                               Tsr29_SPILL_259 <= 64'sh_8000_0000_0000_0000+Tsro29_4_V_1+(rtl_sign_extend4(Tsro29_4_V_0)<<32'sd52);
                               Tsp27_SPILL_256 <= 64'sh1;
                               end 
                              if ((Tsro29_4_V_1==32'sd0/*0:Tsro29.4_V_1*/) && !(32'sd1&(32'sd0/*0:USA36*/==(32'sd512^Tsro29_4_V_6))) && 
                      !Tsfl1_7_V_2)  begin 
                               xpc10 <= 10'sd715/*715:xpc10*/;
                               Tsp27_SPILL_256 <= 64'sh0;
                               Tsro29_4_V_0 <= 16'sh0;
                               end 
                              if ((Tsro29_4_V_1==32'sd0/*0:Tsro29.4_V_1*/) && !(32'sd1&(32'sd0/*0:USA36*/==(32'sd512^Tsro29_4_V_6))) && 
                      Tsfl1_7_V_2)  begin 
                               xpc10 <= 10'sd713/*713:xpc10*/;
                               Tsp27_SPILL_256 <= 64'sh1;
                               Tsro29_4_V_0 <= 16'sh0;
                               end 
                               end 
                      
                  10'sd809/*809:xpc10*/:  begin 
                      if (32'sd1&(32'sd0/*0:USA36*/==(32'sd512^Tsro29_4_V_6)))  begin 
                               xpc10 <= 10'sd810/*810:xpc10*/;
                               Tsro29_4_V_1 <= -64'sh2&Tsro29_4_V_1;
                               end 
                              if (!Tsfl0_9_V_2 && (Tsro29_4_V_1!=32'sd0/*0:Tsro29.4_V_1*/) && !(32'sd1&(32'sd0/*0:USA36*/==(32'sd512^
                      Tsro29_4_V_6))))  begin 
                               xpc10 <= 10'sd812/*812:xpc10*/;
                               Tsr29_SPILL_259 <= Tsro29_4_V_1+(rtl_sign_extend4(Tsro29_4_V_0)<<32'sd52);
                               Tsp27_SPILL_256 <= 64'sh0;
                               end 
                              if (Tsfl0_9_V_2 && (Tsro29_4_V_1!=32'sd0/*0:Tsro29.4_V_1*/) && !(32'sd1&(32'sd0/*0:USA36*/==(32'sd512^Tsro29_4_V_6
                      ))))  begin 
                               xpc10 <= 10'sd812/*812:xpc10*/;
                               Tsr29_SPILL_259 <= 64'sh_8000_0000_0000_0000+Tsro29_4_V_1+(rtl_sign_extend4(Tsro29_4_V_0)<<32'sd52);
                               Tsp27_SPILL_256 <= 64'sh1;
                               end 
                              if (!Tsfl0_9_V_2 && (Tsro29_4_V_1==32'sd0/*0:Tsro29.4_V_1*/) && !(32'sd1&(32'sd0/*0:USA36*/==(32'sd512^
                      Tsro29_4_V_6))))  begin 
                               xpc10 <= 10'sd813/*813:xpc10*/;
                               Tsp27_SPILL_256 <= 64'sh0;
                               Tsro29_4_V_0 <= 16'sh0;
                               end 
                              if (Tsfl0_9_V_2 && (Tsro29_4_V_1==32'sd0/*0:Tsro29.4_V_1*/) && !(32'sd1&(32'sd0/*0:USA36*/==(32'sd512^Tsro29_4_V_6
                      ))))  begin 
                               xpc10 <= 10'sd811/*811:xpc10*/;
                               Tsp27_SPILL_256 <= 64'sh1;
                               Tsro29_4_V_0 <= 16'sh0;
                               end 
                               end 
                      endcase
              if ((Tsco3_7_V_0>=32'sh100_0000)) 
                  case (xpc10)
                      10'sd370/*370:xpc10*/:  begin 
                           xpc10 <= 10'sd374/*374:xpc10*/;
                           Tsco3_7_V_1 <= rtl_unsigned_bitextract3(8'h0+A_8_US_CC_SCALbx14_ARA0[$unsigned((Tsco3_7_V_0>>32'sd24))]);
                           end 
                          
                      10'sd483/*483:xpc10*/:  begin 
                           xpc10 <= 10'sd487/*487:xpc10*/;
                           Tsco3_7_V_1 <= rtl_unsigned_bitextract3(8'h0+A_8_US_CC_SCALbx14_ARA0[$unsigned((Tsco3_7_V_0>>32'sd24))]);
                           end 
                          
                      10'sd494/*494:xpc10*/:  begin 
                           xpc10 <= 10'sd498/*498:xpc10*/;
                           Tsco3_7_V_1 <= rtl_unsigned_bitextract3(8'h0+A_8_US_CC_SCALbx14_ARA0[$unsigned((Tsco3_7_V_0>>32'sd24))]);
                           end 
                          
                      10'sd650/*650:xpc10*/:  begin 
                           xpc10 <= 10'sd654/*654:xpc10*/;
                           Tsco3_7_V_1 <= rtl_unsigned_bitextract3(8'h0+A_8_US_CC_SCALbx14_ARA0[$unsigned((Tsco3_7_V_0>>32'sd24))]);
                           end 
                          
                      10'sd661/*661:xpc10*/:  begin 
                           xpc10 <= 10'sd665/*665:xpc10*/;
                           Tsco3_7_V_1 <= rtl_unsigned_bitextract3(8'h0+A_8_US_CC_SCALbx14_ARA0[$unsigned((Tsco3_7_V_0>>32'sd24))]);
                           end 
                          
                      10'sd748/*748:xpc10*/:  begin 
                           xpc10 <= 10'sd752/*752:xpc10*/;
                           Tsco3_7_V_1 <= rtl_unsigned_bitextract3(8'h0+A_8_US_CC_SCALbx14_ARA0[$unsigned((Tsco3_7_V_0>>32'sd24))]);
                           end 
                          
                      10'sd759/*759:xpc10*/:  begin 
                           xpc10 <= 10'sd763/*763:xpc10*/;
                           Tsco3_7_V_1 <= rtl_unsigned_bitextract3(8'h0+A_8_US_CC_SCALbx14_ARA0[$unsigned((Tsco3_7_V_0>>32'sd24))]);
                           end 
                          endcase
                  
              case (xpc10)
                  10'sd288/*288:xpc10*/:  begin 
                      if (!Tsfl1_22_V_0 && (Tsro28_4_V_1!=32'sd0/*0:Tsro28.4_V_1*/) && !(32'sd1&(32'sd0/*0:USA120*/==(32'sd512^Tsro28_4_V_6
                      ))))  begin 
                               xpc10 <= 10'sd291/*291:xpc10*/;
                               Tsr28_SPILL_259 <= Tsro28_4_V_1+(rtl_sign_extend4(Tsro28_4_V_0)<<32'sd52);
                               Tsp27_SPILL_256 <= 64'sh0;
                               end 
                              if (Tsfl1_22_V_0 && (Tsro28_4_V_1!=32'sd0/*0:Tsro28.4_V_1*/) && !(32'sd1&(32'sd0/*0:USA120*/==(32'sd512
                      ^Tsro28_4_V_6))))  begin 
                               xpc10 <= 10'sd291/*291:xpc10*/;
                               Tsr28_SPILL_259 <= 64'sh_8000_0000_0000_0000+Tsro28_4_V_1+(rtl_sign_extend4(Tsro28_4_V_0)<<32'sd52);
                               Tsp27_SPILL_256 <= 64'sh1;
                               end 
                              if (!Tsfl1_22_V_0 && (Tsro28_4_V_1==32'sd0/*0:Tsro28.4_V_1*/) && !(32'sd1&(32'sd0/*0:USA120*/==(32'sd512
                      ^Tsro28_4_V_6))))  begin 
                               xpc10 <= 10'sd292/*292:xpc10*/;
                               Tsp27_SPILL_256 <= 64'sh0;
                               Tsro28_4_V_0 <= 16'sh0;
                               end 
                              if (Tsfl1_22_V_0 && (Tsro28_4_V_1==32'sd0/*0:Tsro28.4_V_1*/) && !(32'sd1&(32'sd0/*0:USA120*/==(32'sd512
                      ^Tsro28_4_V_6))))  begin 
                               xpc10 <= 10'sd290/*290:xpc10*/;
                               Tsp27_SPILL_256 <= 64'sh1;
                               Tsro28_4_V_0 <= 16'sh0;
                               end 
                              if (32'sd1&(32'sd0/*0:USA120*/==(32'sd512^Tsro28_4_V_6)))  begin 
                               xpc10 <= 10'sd289/*289:xpc10*/;
                               Tsro28_4_V_1 <= -64'sh2&Tsro28_4_V_1;
                               end 
                               end 
                      
                  10'sd810/*810:xpc10*/:  begin 
                      if (!Tsfl0_9_V_2 && (Tsro29_4_V_1!=32'sd0/*0:Tsro29.4_V_1*/))  begin 
                               xpc10 <= 10'sd812/*812:xpc10*/;
                               Tsr29_SPILL_259 <= Tsro29_4_V_1+(rtl_sign_extend4(Tsro29_4_V_0)<<32'sd52);
                               Tsp27_SPILL_256 <= 64'sh0;
                               end 
                              if (Tsfl0_9_V_2 && (Tsro29_4_V_1!=32'sd0/*0:Tsro29.4_V_1*/))  begin 
                               xpc10 <= 10'sd812/*812:xpc10*/;
                               Tsr29_SPILL_259 <= 64'sh_8000_0000_0000_0000+Tsro29_4_V_1+(rtl_sign_extend4(Tsro29_4_V_0)<<32'sd52);
                               Tsp27_SPILL_256 <= 64'sh1;
                               end 
                              if (!Tsfl0_9_V_2 && (Tsro29_4_V_1==32'sd0/*0:Tsro29.4_V_1*/))  begin 
                               xpc10 <= 10'sd813/*813:xpc10*/;
                               Tsp27_SPILL_256 <= 64'sh0;
                               Tsro29_4_V_0 <= 16'sh0;
                               end 
                              if (Tsfl0_9_V_2 && (Tsro29_4_V_1==32'sd0/*0:Tsro29.4_V_1*/))  begin 
                               xpc10 <= 10'sd811/*811:xpc10*/;
                               Tsp27_SPILL_256 <= 64'sh1;
                               Tsro29_4_V_0 <= 16'sh0;
                               end 
                               end 
                      endcase
              if ((32'sd0/*0:USA34*/==(Tsro29_4_V_1<<(32'sd63&rtl_signed_bitextract0(Tsro29_4_V_0))))) 
                  case (xpc10)
                      10'sd717/*717:xpc10*/:  begin 
                           xpc10 <= 10'sd720/*720:xpc10*/;
                           Tss18_SPILL_257 <= Tss18_SPILL_259;
                           Tss18_SPILL_258 <= 64'sh0;
                           end 
                          
                      10'sd815/*815:xpc10*/:  begin 
                           xpc10 <= 10'sd818/*818:xpc10*/;
                           Tss18_SPILL_257 <= Tss18_SPILL_259;
                           Tss18_SPILL_258 <= 64'sh0;
                           end 
                          endcase
                   else 
                  case (xpc10)
                      10'sd717/*717:xpc10*/:  begin 
                           xpc10 <= 10'sd718/*718:xpc10*/;
                           Tss18_SPILL_257 <= Tss18_SPILL_256;
                           Tss18_SPILL_258 <= 64'sh1;
                           end 
                          
                      10'sd815/*815:xpc10*/:  begin 
                           xpc10 <= 10'sd816/*816:xpc10*/;
                           Tss18_SPILL_257 <= Tss18_SPILL_256;
                           Tss18_SPILL_258 <= 64'sh1;
                           end 
                          endcase
              if ((xpc10==10'sd712/*712:xpc10*/))  begin 
                      if ((Tsro29_4_V_1!=32'sd0/*0:Tsro29.4_V_1*/) && !Tsfl1_7_V_2)  begin 
                               xpc10 <= 10'sd714/*714:xpc10*/;
                               Tsr29_SPILL_259 <= Tsro29_4_V_1+(rtl_sign_extend4(Tsro29_4_V_0)<<32'sd52);
                               Tsp27_SPILL_256 <= 64'sh0;
                               end 
                              if ((Tsro29_4_V_1!=32'sd0/*0:Tsro29.4_V_1*/) && Tsfl1_7_V_2)  begin 
                               xpc10 <= 10'sd714/*714:xpc10*/;
                               Tsr29_SPILL_259 <= 64'sh_8000_0000_0000_0000+Tsro29_4_V_1+(rtl_sign_extend4(Tsro29_4_V_0)<<32'sd52);
                               Tsp27_SPILL_256 <= 64'sh1;
                               end 
                              if ((Tsro29_4_V_1==32'sd0/*0:Tsro29.4_V_1*/) && !Tsfl1_7_V_2)  begin 
                               xpc10 <= 10'sd715/*715:xpc10*/;
                               Tsp27_SPILL_256 <= 64'sh0;
                               Tsro29_4_V_0 <= 16'sh0;
                               end 
                              if ((Tsro29_4_V_1==32'sd0/*0:Tsro29.4_V_1*/) && Tsfl1_7_V_2)  begin 
                               xpc10 <= 10'sd713/*713:xpc10*/;
                               Tsp27_SPILL_256 <= 64'sh1;
                               Tsro29_4_V_0 <= 16'sh0;
                               end 
                               end 
                      if (!(!Tsro29_4_V_6)) 
                  case (xpc10)
                      10'sd708/*708:xpc10*/:  xpc10 <= 10'sd709/*709:xpc10*/;

                      10'sd709/*709:xpc10*/:  xpc10 <= 10'sd710/*710:xpc10*/;

                      10'sd806/*806:xpc10*/:  xpc10 <= 10'sd807/*807:xpc10*/;

                      10'sd807/*807:xpc10*/:  xpc10 <= 10'sd808/*808:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      10'sd708/*708:xpc10*/:  begin 
                           xpc10 <= 10'sd711/*711:xpc10*/;
                           Tsro29_4_V_1 <= (Tsro29_4_V_1+rtl_sign_extend4(Tsro29_4_V_5)>>32'sd10);
                           end 
                          
                      10'sd709/*709:xpc10*/:  begin 
                           xpc10 <= 10'sd711/*711:xpc10*/;
                           Tsro29_4_V_1 <= (Tsro29_4_V_1+rtl_sign_extend4(Tsro29_4_V_5)>>32'sd10);
                           end 
                          
                      10'sd806/*806:xpc10*/:  begin 
                           xpc10 <= 10'sd809/*809:xpc10*/;
                           Tsro29_4_V_1 <= (Tsro29_4_V_1+rtl_sign_extend4(Tsro29_4_V_5)>>32'sd10);
                           end 
                          
                      10'sd807/*807:xpc10*/:  begin 
                           xpc10 <= 10'sd809/*809:xpc10*/;
                           Tsro29_4_V_1 <= (Tsro29_4_V_1+rtl_sign_extend4(Tsro29_4_V_5)>>32'sd10);
                           end 
                          endcase
              if (!(!Tsro29_4_V_5)) 
                  case (xpc10)
                      10'sd702/*702:xpc10*/:  begin 
                           xpc10 <= 10'sd705/*705:xpc10*/;
                           Tsr29_SPILL_257 <= Tsr29_SPILL_260;
                           Tsr29_SPILL_258 <= 64'sh0;
                           end 
                          
                      10'sd800/*800:xpc10*/:  begin 
                           xpc10 <= 10'sd803/*803:xpc10*/;
                           Tsr29_SPILL_257 <= Tsr29_SPILL_260;
                           Tsr29_SPILL_258 <= 64'sh0;
                           end 
                          endcase
                   else 
                  case (xpc10)
                      10'sd702/*702:xpc10*/:  begin 
                           xpc10 <= 10'sd703/*703:xpc10*/;
                           Tsr29_SPILL_257 <= Tsr29_SPILL_256;
                           Tsr29_SPILL_258 <= 64'sh1;
                           end 
                          
                      10'sd800/*800:xpc10*/:  begin 
                           xpc10 <= 10'sd801/*801:xpc10*/;
                           Tsr29_SPILL_257 <= Tsr29_SPILL_256;
                           Tsr29_SPILL_258 <= 64'sh1;
                           end 
                          endcase
              if ((Tsmu24_24_V_7<Tsmu24_24_V_5)) 
                  case (xpc10)
                      10'sd688/*688:xpc10*/:  begin 
                           xpc10 <= 10'sd689/*689:xpc10*/;
                           Tsm24_SPILL_262 <= 64'sh1;
                           Tsm24_SPILL_260 <= fastspilldup28;
                           end 
                          
                      10'sd786/*786:xpc10*/:  begin 
                           xpc10 <= 10'sd787/*787:xpc10*/;
                           Tsm24_SPILL_262 <= 64'sh1;
                           Tsm24_SPILL_260 <= fastspilldup18;
                           end 
                          endcase
                   else 
                  case (xpc10)
                      10'sd688/*688:xpc10*/:  begin 
                           xpc10 <= 10'sd725/*725:xpc10*/;
                           Tsm24_SPILL_262 <= 64'sh0;
                           Tsm24_SPILL_260 <= fastspilldup28;
                           end 
                          
                      10'sd786/*786:xpc10*/:  begin 
                           xpc10 <= 10'sd823/*823:xpc10*/;
                           Tsm24_SPILL_262 <= 64'sh0;
                           Tsm24_SPILL_260 <= fastspilldup18;
                           end 
                          endcase
              if ((Tsmu24_24_V_5<Tsmu24_24_V_6)) 
                  case (xpc10)
                      10'sd683/*683:xpc10*/:  begin 
                           xpc10 <= 10'sd684/*684:xpc10*/;
                           Tsm24_SPILL_259 <= 64'sh1;
                           Tsm24_SPILL_257 <= fastspilldup26;
                           end 
                          
                      10'sd781/*781:xpc10*/:  begin 
                           xpc10 <= 10'sd782/*782:xpc10*/;
                           Tsm24_SPILL_259 <= 64'sh1;
                           Tsm24_SPILL_257 <= fastspilldup16;
                           end 
                          endcase
                   else 
                  case (xpc10)
                      10'sd683/*683:xpc10*/:  begin 
                           xpc10 <= 10'sd726/*726:xpc10*/;
                           Tsm24_SPILL_259 <= 64'sh0;
                           Tsm24_SPILL_257 <= fastspilldup26;
                           end 
                          
                      10'sd781/*781:xpc10*/:  begin 
                           xpc10 <= 10'sd824/*824:xpc10*/;
                           Tsm24_SPILL_259 <= 64'sh0;
                           Tsm24_SPILL_257 <= fastspilldup16;
                           end 
                          endcase

              case (xpc10)
                  10'sd289/*289:xpc10*/:  begin 
                      if (!Tsfl1_22_V_0 && (Tsro28_4_V_1!=32'sd0/*0:Tsro28.4_V_1*/))  begin 
                               xpc10 <= 10'sd291/*291:xpc10*/;
                               Tsr28_SPILL_259 <= Tsro28_4_V_1+(rtl_sign_extend4(Tsro28_4_V_0)<<32'sd52);
                               Tsp27_SPILL_256 <= 64'sh0;
                               end 
                              if (Tsfl1_22_V_0 && (Tsro28_4_V_1!=32'sd0/*0:Tsro28.4_V_1*/))  begin 
                               xpc10 <= 10'sd291/*291:xpc10*/;
                               Tsr28_SPILL_259 <= 64'sh_8000_0000_0000_0000+Tsro28_4_V_1+(rtl_sign_extend4(Tsro28_4_V_0)<<32'sd52);
                               Tsp27_SPILL_256 <= 64'sh1;
                               end 
                              if (!Tsfl1_22_V_0 && (Tsro28_4_V_1==32'sd0/*0:Tsro28.4_V_1*/))  begin 
                               xpc10 <= 10'sd292/*292:xpc10*/;
                               Tsp27_SPILL_256 <= 64'sh0;
                               Tsro28_4_V_0 <= 16'sh0;
                               end 
                              if (Tsfl1_22_V_0 && (Tsro28_4_V_1==32'sd0/*0:Tsro28.4_V_1*/))  begin 
                               xpc10 <= 10'sd290/*290:xpc10*/;
                               Tsp27_SPILL_256 <= 64'sh1;
                               Tsro28_4_V_0 <= 16'sh0;
                               end 
                               end 
                      
                  10'sd393/*393:xpc10*/:  begin 
                      if (!Tssu2_4_V_0 && (Tsro0_16_V_1!=32'sd0/*0:Tsro0.16_V_1*/))  begin 
                               xpc10 <= 10'sd395/*395:xpc10*/;
                               Tsr0_SPILL_259 <= Tsro0_16_V_1+(rtl_sign_extend4(Tsro0_16_V_0)<<32'sd52);
                               Tsp27_SPILL_256 <= 64'sh0;
                               end 
                              if (Tssu2_4_V_0 && (Tsro0_16_V_1!=32'sd0/*0:Tsro0.16_V_1*/))  begin 
                               xpc10 <= 10'sd395/*395:xpc10*/;
                               Tsr0_SPILL_259 <= 64'sh_8000_0000_0000_0000+Tsro0_16_V_1+(rtl_sign_extend4(Tsro0_16_V_0)<<32'sd52);
                               Tsp27_SPILL_256 <= 64'sh1;
                               end 
                              if (!Tssu2_4_V_0 && (Tsro0_16_V_1==32'sd0/*0:Tsro0.16_V_1*/))  begin 
                               xpc10 <= 10'sd396/*396:xpc10*/;
                               Tsp27_SPILL_256 <= 64'sh0;
                               Tsro0_16_V_0 <= 16'sh0;
                               end 
                              if (Tssu2_4_V_0 && (Tsro0_16_V_1==32'sd0/*0:Tsro0.16_V_1*/))  begin 
                               xpc10 <= 10'sd394/*394:xpc10*/;
                               Tsp27_SPILL_256 <= 64'sh1;
                               Tsro0_16_V_0 <= 16'sh0;
                               end 
                               end 
                      
                  10'sd551/*551:xpc10*/:  begin 
                      if (!Tsfl1_18_V_2 && (Tsro33_4_V_1!=32'sd0/*0:Tsro33.4_V_1*/))  begin 
                               xpc10 <= 10'sd553/*553:xpc10*/;
                               Tsr33_SPILL_259 <= Tsro33_4_V_1+(rtl_sign_extend4(Tsro33_4_V_0)<<32'sd52);
                               Tsp27_SPILL_256 <= 64'sh0;
                               end 
                              if (Tsfl1_18_V_2 && (Tsro33_4_V_1!=32'sd0/*0:Tsro33.4_V_1*/))  begin 
                               xpc10 <= 10'sd553/*553:xpc10*/;
                               Tsr33_SPILL_259 <= 64'sh_8000_0000_0000_0000+Tsro33_4_V_1+(rtl_sign_extend4(Tsro33_4_V_0)<<32'sd52);
                               Tsp27_SPILL_256 <= 64'sh1;
                               end 
                              if (!Tsfl1_18_V_2 && (Tsro33_4_V_1==32'sd0/*0:Tsro33.4_V_1*/))  begin 
                               xpc10 <= 10'sd554/*554:xpc10*/;
                               Tsp27_SPILL_256 <= 64'sh0;
                               Tsro33_4_V_0 <= 16'sh0;
                               end 
                              if (Tsfl1_18_V_2 && (Tsro33_4_V_1==32'sd0/*0:Tsro33.4_V_1*/))  begin 
                               xpc10 <= 10'sd552/*552:xpc10*/;
                               Tsp27_SPILL_256 <= 64'sh1;
                               Tsro33_4_V_0 <= 16'sh0;
                               end 
                               end 
                      endcase
              if ((32'sd4094/*4094:USA28*/==(64'shfff&(Tspr11_2_V_1>>32'sd51)))) 
                  case (xpc10)
                      10'sd638/*638:xpc10*/:  begin 
                           xpc10 <= 10'sd639/*639:xpc10*/;
                           Tsf0SPILL12_256 <= rtl_sign_extend6((32'sd0/*0:USA32*/==(32'sd0/*0:USA30*/==(64'sh7_ffff_ffff_ffff&Tspr11_2_V_1
                          ))));

                           end 
                          
                      10'sd736/*736:xpc10*/:  begin 
                           xpc10 <= 10'sd737/*737:xpc10*/;
                           Tsf0SPILL12_256 <= rtl_sign_extend6((32'sd0/*0:USA32*/==(32'sd0/*0:USA30*/==(64'sh7_ffff_ffff_ffff&Tspr11_2_V_1
                          ))));

                           end 
                          endcase
                   else 
                  case (xpc10)
                      10'sd638/*638:xpc10*/:  begin 
                           xpc10 <= 10'sd644/*644:xpc10*/;
                           Tspr11_2_V_4 <= 1'h0;
                           Tsf0SPILL12_256 <= 32'sd0;
                           end 
                          
                      10'sd736/*736:xpc10*/:  begin 
                           xpc10 <= 10'sd742/*742:xpc10*/;
                           Tspr11_2_V_4 <= 1'h0;
                           Tsf0SPILL12_256 <= 32'sd0;
                           end 
                          endcase
              if ((32'sd4094/*4094:USA22*/==(64'shfff&(Tspr11_2_V_0>>32'sd51)))) 
                  case (xpc10)
                      10'sd636/*636:xpc10*/:  begin 
                           xpc10 <= 10'sd637/*637:xpc10*/;
                           Tsf0SPILL10_256 <= rtl_sign_extend6((32'sd0/*0:USA26*/==(32'sd0/*0:USA24*/==(64'sh7_ffff_ffff_ffff&Tspr11_2_V_0
                          ))));

                           end 
                          
                      10'sd734/*734:xpc10*/:  begin 
                           xpc10 <= 10'sd735/*735:xpc10*/;
                           Tsf0SPILL10_256 <= rtl_sign_extend6((32'sd0/*0:USA26*/==(32'sd0/*0:USA24*/==(64'sh7_ffff_ffff_ffff&Tspr11_2_V_0
                          ))));

                           end 
                          endcase
                   else 
                  case (xpc10)
                      10'sd636/*636:xpc10*/:  begin 
                           xpc10 <= 10'sd645/*645:xpc10*/;
                           Tspr11_2_V_2 <= 1'h0;
                           Tsf0SPILL10_256 <= 32'sd0;
                           end 
                          
                      10'sd734/*734:xpc10*/:  begin 
                           xpc10 <= 10'sd743/*743:xpc10*/;
                           Tspr11_2_V_2 <= 1'h0;
                           Tsf0SPILL10_256 <= 32'sd0;
                           end 
                          endcase
              if (Tsin1_17_V_0) 
                  case (xpc10)
                      10'sd619/*619:xpc10*/:  begin 
                           xpc10 <= 10'sd620/*620:xpc10*/;
                           Tsi1_SPILL_257 <= -32'sd2*Tdsi3_5_V_2*(32'sd1+32'sd2*Tdsi3_5_V_2);
                           end 
                          
                      10'sd626/*626:xpc10*/:  begin 
                           xpc10 <= 10'sd627/*627:xpc10*/;
                           Tsp5_SPILL_256 <= 64'sh1;
                           Tsin1_17_V_2 <= rtl_unsigned_extend7(Tsin1_17_V_1);
                           end 
                          endcase
                   else 
                  case (xpc10)
                      10'sd619/*619:xpc10*/:  begin 
                           xpc10 <= 10'sd630/*630:xpc10*/;
                           Tsi1_SPILL_257 <= 32'sd2*Tdsi3_5_V_2*(32'sd1+32'sd2*Tdsi3_5_V_2);
                           end 
                          
                      10'sd626/*626:xpc10*/:  begin 
                           xpc10 <= 10'sd629/*629:xpc10*/;
                           Tsp5_SPILL_256 <= 64'sh0;
                           Tsin1_17_V_2 <= rtl_unsigned_extend7(Tsin1_17_V_1);
                           end 
                          endcase
              if (($signed(Tsfl1_18_V_9)<64'sh0)) 
                  case (xpc10)
                      10'sd532/*532:xpc10*/:  begin 
                           xpc10 <= 10'sd564/*564:xpc10*/;
                           Tsfl1_18_V_8 <= -64'd1+Tsfl1_18_V_8;
                           end 
                          
                      10'sd569/*569:xpc10*/:  begin 
                           xpc10 <= 10'sd564/*564:xpc10*/;
                           Tsfl1_18_V_8 <= -64'd1+Tsfl1_18_V_8;
                           end 
                          endcase
                   else 
                  case (xpc10)
                      10'sd532/*532:xpc10*/:  begin 
                           xpc10 <= 10'sd533/*533:xpc10*/;
                           Tsf1SPILL10_260 <= Tsfl1_18_V_8;
                           fastspilldup54 <= Tsfl1_18_V_8;
                           end 
                          
                      10'sd569/*569:xpc10*/:  begin 
                           xpc10 <= 10'sd533/*533:xpc10*/;
                           Tsf1SPILL10_260 <= Tsfl1_18_V_8;
                           fastspilldup54 <= Tsfl1_18_V_8;
                           end 
                          endcase
              if ((xpc10==10'sd259/*259:xpc10*/))  begin 
                      if ((Tsfl0_3_V_0? (64'sh_3ee4_f8b5_88e3_68f1==(64'sh_7fff_ffff_ffff_ffff&Tdsi3_5_V_1)) && Tsfl0_3_V_1: (64'sh_3ee4_f8b5_88e3_68f1
                      ==(64'sh_7fff_ffff_ffff_ffff&Tdsi3_5_V_1)) && !Tsfl0_3_V_1))  begin 
                               xpc10 <= 10'sd263/*263:xpc10*/;
                               Tsf0SPILL14_256 <= 32'sh1;
                               Tsf0SPILL14_258 <= 32'sd1;
                               end 
                              if (Tsfl0_3_V_0 && !Tsfl0_3_V_1)  begin 
                               xpc10 <= 10'sd261/*261:xpc10*/;
                               Tsf0SPILL14_256 <= 32'sh1;
                               Tsf0SPILL14_257 <= 32'sd1;
                               end 
                              if ((Tsfl0_3_V_0? (64'sh_3ee4_f8b5_88e3_68f1!=(64'sh_7fff_ffff_ffff_ffff&Tdsi3_5_V_1)) && Tsfl0_3_V_1: (64'sh_3ee4_f8b5_88e3_68f1
                      !=(64'sh_7fff_ffff_ffff_ffff&Tdsi3_5_V_1)) && !Tsfl0_3_V_1))  begin 
                               xpc10 <= 10'sd262/*262:xpc10*/;
                               Tsf0SPILL14_258 <= $unsigned(Tsfl0_3_V_0^(64'sh_3ee4_f8b5_88e3_68f1<$signed(64'sh_7fff_ffff_ffff_ffff&
                              Tdsi3_5_V_1)));

                               end 
                              if (!Tsfl0_3_V_0 && Tsfl0_3_V_1)  begin 
                               xpc10 <= 10'sd260/*260:xpc10*/;
                               Tsf0SPILL14_257 <= rtl_sign_extend6((32'sd0/*0:USA170*/==((64'sh_3ee4_f8b5_88e3_68f1|64'sh_7fff_ffff_ffff_ffff
                              &Tdsi3_5_V_1)<<32'sd1)));

                               end 
                               end 
                      if ((32'sd4094/*4094:USA16*/==(64'shfff&(Tspr4_3_V_1>>32'sd51)))) 
                  case (xpc10)
                      10'sd188/*188:xpc10*/:  begin 
                           xpc10 <= 10'sd189/*189:xpc10*/;
                           Tsf0SPILL12_256 <= rtl_sign_extend6((32'sd0/*0:USA20*/==(32'sd0/*0:USA18*/==(64'sh7_ffff_ffff_ffff&Tspr4_3_V_1
                          ))));

                           end 
                          
                      10'sd206/*206:xpc10*/:  begin 
                           xpc10 <= 10'sd207/*207:xpc10*/;
                           Tsf0SPILL12_256 <= rtl_sign_extend6((32'sd0/*0:USA20*/==(32'sd0/*0:USA18*/==(64'sh7_ffff_ffff_ffff&Tspr4_3_V_1
                          ))));

                           end 
                          endcase
                   else 
                  case (xpc10)
                      10'sd188/*188:xpc10*/:  begin 
                           xpc10 <= 10'sd729/*729:xpc10*/;
                           Tspr4_3_V_4 <= 1'h0;
                           Tsf0SPILL12_256 <= 32'sd0;
                           end 
                          
                      10'sd206/*206:xpc10*/:  begin 
                           xpc10 <= 10'sd631/*631:xpc10*/;
                           Tspr4_3_V_4 <= 1'h0;
                           Tsf0SPILL12_256 <= 32'sd0;
                           end 
                          endcase
              if ((32'sd4094/*4094:USA10*/==(64'shfff&(Tspr4_3_V_0>>32'sd51)))) 
                  case (xpc10)
                      10'sd186/*186:xpc10*/:  begin 
                           xpc10 <= 10'sd187/*187:xpc10*/;
                           Tsf0SPILL10_256 <= rtl_sign_extend6((32'sd0/*0:USA14*/==(32'sd0/*0:USA12*/==(64'sh7_ffff_ffff_ffff&Tspr4_3_V_0
                          ))));

                           end 
                          
                      10'sd204/*204:xpc10*/:  begin 
                           xpc10 <= 10'sd205/*205:xpc10*/;
                           Tsf0SPILL10_256 <= rtl_sign_extend6((32'sd0/*0:USA14*/==(32'sd0/*0:USA12*/==(64'sh7_ffff_ffff_ffff&Tspr4_3_V_0
                          ))));

                           end 
                          endcase
                   else 
                  case (xpc10)
                      10'sd186/*186:xpc10*/:  begin 
                           xpc10 <= 10'sd730/*730:xpc10*/;
                           Tspr4_3_V_2 <= 1'h0;
                           Tsf0SPILL10_256 <= 32'sd0;
                           end 
                          
                      10'sd204/*204:xpc10*/:  begin 
                           xpc10 <= 10'sd632/*632:xpc10*/;
                           Tspr4_3_V_2 <= 1'h0;
                           Tsf0SPILL10_256 <= 32'sd0;
                           end 
                          endcase

              case (xpc10)
                  10'sd267/*267:xpc10*/:  begin 
                      if (!(!(!rtl_signed_bitextract0(Tsad1_3_V_6))))  begin 
                               xpc10 <= 10'sd268/*268:xpc10*/;
                               Tsad1_3_V_4 <= Tsad1_3_V_4;
                               Tssh8_5_V_0 <= Tsad1_3_V_4;
                               end 
                              if (!(!rtl_signed_bitextract0(Tsad1_3_V_6)) && (rtl_signed_bitextract0(Tsad1_3_V_6)>=32'sd64) && (Tsad1_3_V_4
                      ==32'sd0/*0:Tsad1.3_V_4*/))  begin 
                               xpc10 <= 10'sd307/*307:xpc10*/;
                               Tssh8_5_V_0 <= 64'h0;
                               end 
                              if (!(!rtl_signed_bitextract0(Tsad1_3_V_6)) && (rtl_signed_bitextract0(Tsad1_3_V_6)>=32'sd64) && (Tsad1_3_V_4
                      !=32'sd0/*0:Tsad1.3_V_4*/))  begin 
                               xpc10 <= 10'sd307/*307:xpc10*/;
                               Tssh8_5_V_0 <= 64'h1;
                               end 
                              if (!(!rtl_signed_bitextract0(Tsad1_3_V_6)) && (rtl_signed_bitextract0(Tsad1_3_V_6)<32'sd64))  begin 
                               xpc10 <= 10'sd301/*301:xpc10*/;
                               fastspilldup60 <= (Tsad1_3_V_4>>(32'sd63&rtl_signed_bitextract0(Tsad1_3_V_6)));
                               end 
                               end 
                      
                  10'sd308/*308:xpc10*/:  begin 
                      if (!(!(!rtl_signed_bitextract0(Tsad1_3_V_6))))  begin 
                               xpc10 <= 10'sd268/*268:xpc10*/;
                               Tsad1_3_V_4 <= Tsad1_3_V_4;
                               Tssh8_5_V_0 <= Tsad1_3_V_4;
                               end 
                              if (!(!rtl_signed_bitextract0(Tsad1_3_V_6)) && (rtl_signed_bitextract0(Tsad1_3_V_6)>=32'sd64) && (Tsad1_3_V_4
                      ==32'sd0/*0:Tsad1.3_V_4*/))  begin 
                               xpc10 <= 10'sd307/*307:xpc10*/;
                               Tssh8_5_V_0 <= 64'h0;
                               end 
                              if (!(!rtl_signed_bitextract0(Tsad1_3_V_6)) && (rtl_signed_bitextract0(Tsad1_3_V_6)>=32'sd64) && (Tsad1_3_V_4
                      !=32'sd0/*0:Tsad1.3_V_4*/))  begin 
                               xpc10 <= 10'sd307/*307:xpc10*/;
                               Tssh8_5_V_0 <= 64'h1;
                               end 
                              if (!(!rtl_signed_bitextract0(Tsad1_3_V_6)) && (rtl_signed_bitextract0(Tsad1_3_V_6)<32'sd64))  begin 
                               xpc10 <= 10'sd301/*301:xpc10*/;
                               fastspilldup60 <= (Tsad1_3_V_4>>(32'sd63&rtl_signed_bitextract0(Tsad1_3_V_6)));
                               end 
                               end 
                      
                  10'sd320/*320:xpc10*/:  begin 
                      if (!(!(!rtl_signed_bitextract0((0-Tsad1_3_V_6)))))  begin 
                               xpc10 <= 10'sd321/*321:xpc10*/;
                               Tsad1_3_V_3 <= Tsad1_3_V_3;
                               Tssh17_6_V_0 <= Tsad1_3_V_3;
                               end 
                              if ((Tsad1_3_V_3==32'sd0/*0:Tsad1.3_V_3*/) && !(!rtl_signed_bitextract0((0-Tsad1_3_V_6))) && (rtl_signed_bitextract0((0
                      -Tsad1_3_V_6))>=32'sd64))  begin 
                               xpc10 <= 10'sd328/*328:xpc10*/;
                               Tssh17_6_V_0 <= 64'h0;
                               end 
                              if ((Tsad1_3_V_3!=32'sd0/*0:Tsad1.3_V_3*/) && !(!rtl_signed_bitextract0((0-Tsad1_3_V_6))) && (rtl_signed_bitextract0((0
                      -Tsad1_3_V_6))>=32'sd64))  begin 
                               xpc10 <= 10'sd328/*328:xpc10*/;
                               Tssh17_6_V_0 <= 64'h1;
                               end 
                              if (!(!rtl_signed_bitextract0((0-Tsad1_3_V_6))) && (rtl_signed_bitextract0((0-Tsad1_3_V_6))<32'sd64))  begin 
                               xpc10 <= 10'sd322/*322:xpc10*/;
                               fastspilldup62 <= (Tsad1_3_V_3>>(32'sd63&rtl_signed_bitextract0((0-Tsad1_3_V_6))));
                               end 
                               end 
                      
                  10'sd329/*329:xpc10*/:  begin 
                      if (!(!(!rtl_signed_bitextract0((0-Tsad1_3_V_6)))))  begin 
                               xpc10 <= 10'sd321/*321:xpc10*/;
                               Tsad1_3_V_3 <= Tsad1_3_V_3;
                               Tssh17_6_V_0 <= Tsad1_3_V_3;
                               end 
                              if ((Tsad1_3_V_3==32'sd0/*0:Tsad1.3_V_3*/) && !(!rtl_signed_bitextract0((0-Tsad1_3_V_6))) && (rtl_signed_bitextract0((0
                      -Tsad1_3_V_6))>=32'sd64))  begin 
                               xpc10 <= 10'sd328/*328:xpc10*/;
                               Tssh17_6_V_0 <= 64'h0;
                               end 
                              if ((Tsad1_3_V_3!=32'sd0/*0:Tsad1.3_V_3*/) && !(!rtl_signed_bitextract0((0-Tsad1_3_V_6))) && (rtl_signed_bitextract0((0
                      -Tsad1_3_V_6))>=32'sd64))  begin 
                               xpc10 <= 10'sd328/*328:xpc10*/;
                               Tssh17_6_V_0 <= 64'h1;
                               end 
                              if (!(!rtl_signed_bitextract0((0-Tsad1_3_V_6))) && (rtl_signed_bitextract0((0-Tsad1_3_V_6))<32'sd64))  begin 
                               xpc10 <= 10'sd322/*322:xpc10*/;
                               fastspilldup62 <= (Tsad1_3_V_3>>(32'sd63&rtl_signed_bitextract0((0-Tsad1_3_V_6))));
                               end 
                               end 
                      
                  10'sd364/*364:xpc10*/:  begin 
                      if (!(!(!rtl_signed_bitextract0(Tssu2_4_V_7))))  begin 
                               xpc10 <= 10'sd365/*365:xpc10*/;
                               Tssu2_4_V_5 <= Tssu2_4_V_5;
                               Tssh32_5_V_0 <= Tssu2_4_V_5;
                               end 
                              if (!(!rtl_signed_bitextract0(Tssu2_4_V_7)) && (rtl_signed_bitextract0(Tssu2_4_V_7)>=32'sd64) && (Tssu2_4_V_5
                      ==32'sd0/*0:Tssu2.4_V_5*/))  begin 
                               xpc10 <= 10'sd411/*411:xpc10*/;
                               Tssh32_5_V_0 <= 64'h0;
                               end 
                              if (!(!rtl_signed_bitextract0(Tssu2_4_V_7)) && (rtl_signed_bitextract0(Tssu2_4_V_7)>=32'sd64) && (Tssu2_4_V_5
                      !=32'sd0/*0:Tssu2.4_V_5*/))  begin 
                               xpc10 <= 10'sd411/*411:xpc10*/;
                               Tssh32_5_V_0 <= 64'h1;
                               end 
                              if (!(!rtl_signed_bitextract0(Tssu2_4_V_7)) && (rtl_signed_bitextract0(Tssu2_4_V_7)<32'sd64))  begin 
                               xpc10 <= 10'sd406/*406:xpc10*/;
                               fastspilldup70 <= (Tssu2_4_V_5>>(32'sd63&rtl_signed_bitextract0(Tssu2_4_V_7)));
                               end 
                               end 
                      
                  10'sd412/*412:xpc10*/:  begin 
                      if (!(!(!rtl_signed_bitextract0(Tssu2_4_V_7))))  begin 
                               xpc10 <= 10'sd365/*365:xpc10*/;
                               Tssu2_4_V_5 <= Tssu2_4_V_5;
                               Tssh32_5_V_0 <= Tssu2_4_V_5;
                               end 
                              if (!(!rtl_signed_bitextract0(Tssu2_4_V_7)) && (rtl_signed_bitextract0(Tssu2_4_V_7)>=32'sd64) && (Tssu2_4_V_5
                      ==32'sd0/*0:Tssu2.4_V_5*/))  begin 
                               xpc10 <= 10'sd411/*411:xpc10*/;
                               Tssh32_5_V_0 <= 64'h0;
                               end 
                              if (!(!rtl_signed_bitextract0(Tssu2_4_V_7)) && (rtl_signed_bitextract0(Tssu2_4_V_7)>=32'sd64) && (Tssu2_4_V_5
                      !=32'sd0/*0:Tssu2.4_V_5*/))  begin 
                               xpc10 <= 10'sd411/*411:xpc10*/;
                               Tssh32_5_V_0 <= 64'h1;
                               end 
                              if (!(!rtl_signed_bitextract0(Tssu2_4_V_7)) && (rtl_signed_bitextract0(Tssu2_4_V_7)<32'sd64))  begin 
                               xpc10 <= 10'sd406/*406:xpc10*/;
                               fastspilldup70 <= (Tssu2_4_V_5>>(32'sd63&rtl_signed_bitextract0(Tssu2_4_V_7)));
                               end 
                               end 
                      
                  10'sd424/*424:xpc10*/:  begin 
                      if (!(!(!rtl_signed_bitextract0((0-Tssu2_4_V_7)))))  begin 
                               xpc10 <= 10'sd425/*425:xpc10*/;
                               Tssu2_4_V_4 <= Tssu2_4_V_4;
                               Tssh23_6_V_0 <= Tssu2_4_V_4;
                               end 
                              if ((Tssu2_4_V_4==32'sd0/*0:Tssu2.4_V_4*/) && !(!rtl_signed_bitextract0((0-Tssu2_4_V_7))) && (rtl_signed_bitextract0((0
                      -Tssu2_4_V_7))>=32'sd64))  begin 
                               xpc10 <= 10'sd434/*434:xpc10*/;
                               Tssh23_6_V_0 <= 64'h0;
                               end 
                              if ((Tssu2_4_V_4!=32'sd0/*0:Tssu2.4_V_4*/) && !(!rtl_signed_bitextract0((0-Tssu2_4_V_7))) && (rtl_signed_bitextract0((0
                      -Tssu2_4_V_7))>=32'sd64))  begin 
                               xpc10 <= 10'sd434/*434:xpc10*/;
                               Tssh23_6_V_0 <= 64'h1;
                               end 
                              if (!(!rtl_signed_bitextract0((0-Tssu2_4_V_7))) && (rtl_signed_bitextract0((0-Tssu2_4_V_7))<32'sd64))  begin 
                               xpc10 <= 10'sd429/*429:xpc10*/;
                               fastspilldup68 <= (Tssu2_4_V_4>>(32'sd63&rtl_signed_bitextract0((0-Tssu2_4_V_7))));
                               end 
                               end 
                      
                  10'sd435/*435:xpc10*/:  begin 
                      if (!(!(!rtl_signed_bitextract0((0-Tssu2_4_V_7)))))  begin 
                               xpc10 <= 10'sd425/*425:xpc10*/;
                               Tssu2_4_V_4 <= Tssu2_4_V_4;
                               Tssh23_6_V_0 <= Tssu2_4_V_4;
                               end 
                              if ((Tssu2_4_V_4==32'sd0/*0:Tssu2.4_V_4*/) && !(!rtl_signed_bitextract0((0-Tssu2_4_V_7))) && (rtl_signed_bitextract0((0
                      -Tssu2_4_V_7))>=32'sd64))  begin 
                               xpc10 <= 10'sd434/*434:xpc10*/;
                               Tssh23_6_V_0 <= 64'h0;
                               end 
                              if ((Tssu2_4_V_4!=32'sd0/*0:Tssu2.4_V_4*/) && !(!rtl_signed_bitextract0((0-Tssu2_4_V_7))) && (rtl_signed_bitextract0((0
                      -Tssu2_4_V_7))>=32'sd64))  begin 
                               xpc10 <= 10'sd434/*434:xpc10*/;
                               Tssh23_6_V_0 <= 64'h1;
                               end 
                              if (!(!rtl_signed_bitextract0((0-Tssu2_4_V_7))) && (rtl_signed_bitextract0((0-Tssu2_4_V_7))<32'sd64))  begin 
                               xpc10 <= 10'sd429/*429:xpc10*/;
                               fastspilldup68 <= (Tssu2_4_V_4>>(32'sd63&rtl_signed_bitextract0((0-Tssu2_4_V_7))));
                               end 
                               end 
                      
                  10'sd491/*491:xpc10*/:  begin 
                      if ((Tsfl1_18_V_6!=32'sd0/*0:Tsfl1.18_V_6*/) && !Tsfl1_18_V_3)  begin 
                               xpc10 <= 10'sd493/*493:xpc10*/;
                               Tsco0_2_V_1 <= 8'h0;
                               Tsco0_2_V_0 <= Tsfl1_18_V_6;
                               end 
                              if (!(!Tsfl1_18_V_3))  begin 
                               xpc10 <= 10'sd503/*503:xpc10*/;
                               Tsfl1_18_V_5 <= rtl_signed_bitextract0(rtl_sign_extend2(16'sd1021)+rtl_sign_extend2(Tsfl1_18_V_3)+(0-Tsfl1_18_V_4
                              ));

                               end 
                              if ((Tsfl1_18_V_6==32'sd0/*0:Tsfl1.18_V_6*/) && !Tsfl1_18_V_2 && !Tsfl1_18_V_3)  begin 
                               xpc10 <= 10'sd492/*492:xpc10*/;
                               Tsf1SPILL10_256 <= 64'h0;
                               end 
                              if ((Tsfl1_18_V_6==32'sd0/*0:Tsfl1.18_V_6*/) && Tsfl1_18_V_2 && !Tsfl1_18_V_3)  begin 
                               xpc10 <= 10'sd492/*492:xpc10*/;
                               Tsf1SPILL10_256 <= 64'h_8000_0000_0000_0000;
                               end 
                               end 
                      
                  10'sd642/*642:xpc10*/:  begin 
                      if (!Tspr11_2_V_2 && !Tspr11_2_V_4 && !Tspr11_2_V_3)  begin 
                               xpc10 <= 10'sd643/*643:xpc10*/;
                               Tsf1_SPILL_256 <= Tspr11_2_V_0;
                               end 
                              if (!Tspr11_2_V_2 && !Tspr11_2_V_4 && Tspr11_2_V_3)  begin 
                               xpc10 <= 10'sd643/*643:xpc10*/;
                               Tsf1_SPILL_256 <= Tspr11_2_V_1;
                               end 
                              if (Tspr11_2_V_2 && !Tspr11_2_V_4)  begin 
                               xpc10 <= 10'sd643/*643:xpc10*/;
                               Tsf1_SPILL_256 <= Tspr11_2_V_0;
                               end 
                              if (Tspr11_2_V_4)  begin 
                               xpc10 <= 10'sd643/*643:xpc10*/;
                               Tsf1_SPILL_256 <= Tspr11_2_V_1;
                               end 
                               end 
                      
                  10'sd658/*658:xpc10*/:  begin 
                      if ((Tsfl1_7_V_7!=32'sd0/*0:Tsfl1.7_V_7*/) && !Tsfl1_7_V_4)  begin 
                               xpc10 <= 10'sd660/*660:xpc10*/;
                               Tsco0_2_V_1 <= 8'h0;
                               Tsco0_2_V_0 <= Tsfl1_7_V_7;
                               end 
                              if (!(!Tsfl1_7_V_4))  begin 
                               xpc10 <= 10'sd670/*670:xpc10*/;
                               Tsfl1_7_V_5 <= rtl_signed_bitextract0(-16'sd1023+Tsfl1_7_V_3+Tsfl1_7_V_4);
                               end 
                              if ((Tsfl1_7_V_7==32'sd0/*0:Tsfl1.7_V_7*/) && !Tsfl1_7_V_4 && !Tsfl1_7_V_2)  begin 
                               xpc10 <= 10'sd659/*659:xpc10*/;
                               Tsf1_SPILL_256 <= 64'h0;
                               end 
                              if ((Tsfl1_7_V_7==32'sd0/*0:Tsfl1.7_V_7*/) && !Tsfl1_7_V_4 && Tsfl1_7_V_2)  begin 
                               xpc10 <= 10'sd659/*659:xpc10*/;
                               Tsf1_SPILL_256 <= 64'h_8000_0000_0000_0000;
                               end 
                               end 
                      
                  10'sd740/*740:xpc10*/:  begin 
                      if (!Tspr11_2_V_2 && !Tspr11_2_V_4 && !Tspr11_2_V_3)  begin 
                               xpc10 <= 10'sd741/*741:xpc10*/;
                               Tsf0_SPILL_256 <= Tspr11_2_V_0;
                               end 
                              if (!Tspr11_2_V_2 && !Tspr11_2_V_4 && Tspr11_2_V_3)  begin 
                               xpc10 <= 10'sd741/*741:xpc10*/;
                               Tsf0_SPILL_256 <= Tspr11_2_V_1;
                               end 
                              if (Tspr11_2_V_2 && !Tspr11_2_V_4)  begin 
                               xpc10 <= 10'sd741/*741:xpc10*/;
                               Tsf0_SPILL_256 <= Tspr11_2_V_0;
                               end 
                              if (Tspr11_2_V_4)  begin 
                               xpc10 <= 10'sd741/*741:xpc10*/;
                               Tsf0_SPILL_256 <= Tspr11_2_V_1;
                               end 
                               end 
                      
                  10'sd756/*756:xpc10*/:  begin 
                      if ((Tsfl0_9_V_7!=32'sd0/*0:Tsfl0.9_V_7*/) && !Tsfl0_9_V_4)  begin 
                               xpc10 <= 10'sd758/*758:xpc10*/;
                               Tsco0_2_V_1 <= 8'h0;
                               Tsco0_2_V_0 <= Tsfl0_9_V_7;
                               end 
                              if (!(!Tsfl0_9_V_4))  begin 
                               xpc10 <= 10'sd768/*768:xpc10*/;
                               Tsfl0_9_V_5 <= rtl_signed_bitextract0(-16'sd1023+Tsfl0_9_V_3+Tsfl0_9_V_4);
                               end 
                              if ((Tsfl0_9_V_7==32'sd0/*0:Tsfl0.9_V_7*/) && !Tsfl0_9_V_4 && !Tsfl0_9_V_2)  begin 
                               xpc10 <= 10'sd757/*757:xpc10*/;
                               Tsf0_SPILL_256 <= 64'h0;
                               end 
                              if ((Tsfl0_9_V_7==32'sd0/*0:Tsfl0.9_V_7*/) && !Tsfl0_9_V_4 && Tsfl0_9_V_2)  begin 
                               xpc10 <= 10'sd757/*757:xpc10*/;
                               Tsf0_SPILL_256 <= 64'h_8000_0000_0000_0000;
                               end 
                               end 
                      endcase
              if (!Tspr11_2_V_2 && !Tspr11_2_V_4 && !Tspr11_2_V_3) 
                  case (xpc10)
                      10'sd641/*641:xpc10*/:  begin 
                           xpc10 <= 10'sd643/*643:xpc10*/;
                           Tsf1_SPILL_256 <= Tspr11_2_V_0;
                           end 
                          
                      10'sd739/*739:xpc10*/:  begin 
                           xpc10 <= 10'sd741/*741:xpc10*/;
                           Tsf0_SPILL_256 <= Tspr11_2_V_0;
                           end 
                          endcase
                  if (!Tspr11_2_V_2 && !Tspr11_2_V_4 && Tspr11_2_V_3) 
                  case (xpc10)
                      10'sd641/*641:xpc10*/:  begin 
                           xpc10 <= 10'sd643/*643:xpc10*/;
                           Tsf1_SPILL_256 <= Tspr11_2_V_1;
                           end 
                          
                      10'sd739/*739:xpc10*/:  begin 
                           xpc10 <= 10'sd741/*741:xpc10*/;
                           Tsf0_SPILL_256 <= Tspr11_2_V_1;
                           end 
                          endcase
                  if ((xpc10==10'sd621/*621:xpc10*/))  begin 
                      if ((Tsco5_4_V_0>=32'sh1_0000) && (Tsco5_4_V_0<32'sh100_0000))  begin 
                               xpc10 <= 10'sd624/*624:xpc10*/;
                               Tsco5_4_V_0 <= (Tsco5_4_V_0<<32'sd8);
                               Tsco5_4_V_1 <= 8'h8;
                               end 
                              if ((Tsco5_4_V_0<32'sh1_0000))  begin 
                               xpc10 <= 10'sd622/*622:xpc10*/;
                               Tsco5_4_V_0 <= (Tsco5_4_V_0<<32'sd16);
                               Tsco5_4_V_1 <= 8'h10;
                               end 
                              if ((Tsco5_4_V_0>=32'sh100_0000))  begin 
                               xpc10 <= 10'sd625/*625:xpc10*/;
                               Tsco5_4_V_1 <= rtl_unsigned_bitextract3(8'h0+A_8_US_CC_SCALbx14_ARA0[$unsigned((Tsco5_4_V_0>>32'sd24))]
                              );

                               end 
                               end 
                      if (($signed(Tses25_5_V_2)<64'sh0)) 
                  case (xpc10)
                      10'sd599/*599:xpc10*/:  begin 
                           xpc10 <= 10'sd605/*605:xpc10*/;
                           Tses25_5_V_6 <= -64'sh1_0000_0000+Tses25_5_V_6;
                           end 
                          
                      10'sd611/*611:xpc10*/:  begin 
                           xpc10 <= 10'sd605/*605:xpc10*/;
                           Tses25_5_V_6 <= -64'sh1_0000_0000+Tses25_5_V_6;
                           end 
                          endcase
                   else 
                  case (xpc10)
                      10'sd599/*599:xpc10*/:  begin 
                           xpc10 <= 10'sd600/*600:xpc10*/;
                           Tses25_5_V_2 <= (Tses25_5_V_2<<32'sd32)|(Tses25_5_V_3>>32'sd32);
                           end 
                          
                      10'sd611/*611:xpc10*/:  begin 
                           xpc10 <= 10'sd600/*600:xpc10*/;
                           Tses25_5_V_2 <= (Tses25_5_V_2<<32'sd32)|(Tses25_5_V_3>>32'sd32);
                           end 
                          endcase
              if (Tsfl1_18_V_2) 
                  case (xpc10)
                      10'sd480/*480:xpc10*/:  begin 
                           xpc10 <= 10'sd481/*481:xpc10*/;
                           Tsf1SPILL10_256 <= 64'h_fff0_0000_0000_0000;
                           end 
                          
                      10'sd539/*539:xpc10*/:  begin 
                           xpc10 <= 10'sd540/*540:xpc10*/;
                           fastspilldup56 <= 64'h_fff0_0000_0000_0000;
                           end 
                          endcase
                   else 
                  case (xpc10)
                      10'sd480/*480:xpc10*/:  begin 
                           xpc10 <= 10'sd481/*481:xpc10*/;
                           Tsf1SPILL10_256 <= 64'h_7ff0_0000_0000_0000;
                           end 
                          
                      10'sd539/*539:xpc10*/:  begin 
                           xpc10 <= 10'sd540/*540:xpc10*/;
                           fastspilldup56 <= 64'h_7ff0_0000_0000_0000;
                           end 
                          endcase

              case (xpc10)
                  10'sd315/*315:xpc10*/:  begin 
                      if (!Tspr12_2_V_2 && !Tspr12_2_V_4 && !Tspr12_2_V_3)  begin 
                               xpc10 <= 10'sd316/*316:xpc10*/;
                               Tsa1_SPILL_256 <= Tspr12_2_V_0;
                               end 
                              if (!Tspr12_2_V_2 && !Tspr12_2_V_4 && Tspr12_2_V_3)  begin 
                               xpc10 <= 10'sd316/*316:xpc10*/;
                               Tsa1_SPILL_256 <= Tspr12_2_V_1;
                               end 
                              if (Tspr12_2_V_2 && !Tspr12_2_V_4)  begin 
                               xpc10 <= 10'sd316/*316:xpc10*/;
                               Tsa1_SPILL_256 <= Tspr12_2_V_0;
                               end 
                              if (Tspr12_2_V_4)  begin 
                               xpc10 <= 10'sd316/*316:xpc10*/;
                               Tsa1_SPILL_256 <= Tspr12_2_V_1;
                               end 
                               end 
                      
                  10'sd336/*336:xpc10*/:  begin 
                      if (!Tspr21_3_V_2 && !Tspr21_3_V_4 && !Tspr21_3_V_3)  begin 
                               xpc10 <= 10'sd337/*337:xpc10*/;
                               Tsa1_SPILL_256 <= Tspr21_3_V_0;
                               end 
                              if (!Tspr21_3_V_2 && !Tspr21_3_V_4 && Tspr21_3_V_3)  begin 
                               xpc10 <= 10'sd337/*337:xpc10*/;
                               Tsa1_SPILL_256 <= Tspr21_3_V_1;
                               end 
                              if (Tspr21_3_V_2 && !Tspr21_3_V_4)  begin 
                               xpc10 <= 10'sd337/*337:xpc10*/;
                               Tsa1_SPILL_256 <= Tspr21_3_V_0;
                               end 
                              if (Tspr21_3_V_4)  begin 
                               xpc10 <= 10'sd337/*337:xpc10*/;
                               Tsa1_SPILL_256 <= Tspr21_3_V_1;
                               end 
                               end 
                      
                  10'sd359/*359:xpc10*/:  begin 
                      if (!Tspr27_2_V_2 && !Tspr27_2_V_4 && !Tspr27_2_V_3)  begin 
                               xpc10 <= 10'sd360/*360:xpc10*/;
                               Tss2_SPILL_256 <= Tspr27_2_V_0;
                               end 
                              if (!Tspr27_2_V_2 && !Tspr27_2_V_4 && Tspr27_2_V_3)  begin 
                               xpc10 <= 10'sd360/*360:xpc10*/;
                               Tss2_SPILL_256 <= Tspr27_2_V_1;
                               end 
                              if (Tspr27_2_V_2 && !Tspr27_2_V_4)  begin 
                               xpc10 <= 10'sd360/*360:xpc10*/;
                               Tss2_SPILL_256 <= Tspr27_2_V_0;
                               end 
                              if (Tspr27_2_V_4)  begin 
                               xpc10 <= 10'sd360/*360:xpc10*/;
                               Tss2_SPILL_256 <= Tspr27_2_V_1;
                               end 
                               end 
                      
                  10'sd419/*419:xpc10*/:  begin 
                      if (!Tspr18_2_V_2 && !Tspr18_2_V_4 && !Tspr18_2_V_3)  begin 
                               xpc10 <= 10'sd420/*420:xpc10*/;
                               Tss2_SPILL_256 <= Tspr18_2_V_0;
                               end 
                              if (!Tspr18_2_V_2 && !Tspr18_2_V_4 && Tspr18_2_V_3)  begin 
                               xpc10 <= 10'sd420/*420:xpc10*/;
                               Tss2_SPILL_256 <= Tspr18_2_V_1;
                               end 
                              if (Tspr18_2_V_2 && !Tspr18_2_V_4)  begin 
                               xpc10 <= 10'sd420/*420:xpc10*/;
                               Tss2_SPILL_256 <= Tspr18_2_V_0;
                               end 
                              if (Tspr18_2_V_4)  begin 
                               xpc10 <= 10'sd420/*420:xpc10*/;
                               Tss2_SPILL_256 <= Tspr18_2_V_1;
                               end 
                               end 
                      
                  10'sd442/*442:xpc10*/:  begin 
                      if (!Tspr7_3_V_2 && !Tspr7_3_V_4 && !Tspr7_3_V_3)  begin 
                               xpc10 <= 10'sd443/*443:xpc10*/;
                               Tss2_SPILL_256 <= Tspr7_3_V_0;
                               end 
                              if (!Tspr7_3_V_2 && !Tspr7_3_V_4 && Tspr7_3_V_3)  begin 
                               xpc10 <= 10'sd443/*443:xpc10*/;
                               Tss2_SPILL_256 <= Tspr7_3_V_1;
                               end 
                              if (Tspr7_3_V_2 && !Tspr7_3_V_4)  begin 
                               xpc10 <= 10'sd443/*443:xpc10*/;
                               Tss2_SPILL_256 <= Tspr7_3_V_0;
                               end 
                              if (Tspr7_3_V_4)  begin 
                               xpc10 <= 10'sd443/*443:xpc10*/;
                               Tss2_SPILL_256 <= Tspr7_3_V_1;
                               end 
                               end 
                      
                  10'sd459/*459:xpc10*/:  begin 
                      if (!Tspr5_2_V_2 && !Tspr5_2_V_4 && !Tspr5_2_V_3)  begin 
                               xpc10 <= 10'sd460/*460:xpc10*/;
                               Tsf1SPILL10_256 <= Tspr5_2_V_0;
                               end 
                              if (!Tspr5_2_V_2 && !Tspr5_2_V_4 && Tspr5_2_V_3)  begin 
                               xpc10 <= 10'sd460/*460:xpc10*/;
                               Tsf1SPILL10_256 <= Tspr5_2_V_1;
                               end 
                              if (Tspr5_2_V_2 && !Tspr5_2_V_4)  begin 
                               xpc10 <= 10'sd460/*460:xpc10*/;
                               Tsf1SPILL10_256 <= Tspr5_2_V_0;
                               end 
                              if (Tspr5_2_V_4)  begin 
                               xpc10 <= 10'sd460/*460:xpc10*/;
                               Tsf1SPILL10_256 <= Tspr5_2_V_1;
                               end 
                               end 
                      
                  10'sd474/*474:xpc10*/:  begin 
                      if (!Tspr10_2_V_2 && !Tspr10_2_V_4 && !Tspr10_2_V_3)  begin 
                               xpc10 <= 10'sd475/*475:xpc10*/;
                               Tsf1SPILL10_256 <= Tspr10_2_V_0;
                               end 
                              if (!Tspr10_2_V_2 && !Tspr10_2_V_4 && Tspr10_2_V_3)  begin 
                               xpc10 <= 10'sd475/*475:xpc10*/;
                               Tsf1SPILL10_256 <= Tspr10_2_V_1;
                               end 
                              if (Tspr10_2_V_2 && !Tspr10_2_V_4)  begin 
                               xpc10 <= 10'sd475/*475:xpc10*/;
                               Tsf1SPILL10_256 <= Tspr10_2_V_0;
                               end 
                              if (Tspr10_2_V_4)  begin 
                               xpc10 <= 10'sd475/*475:xpc10*/;
                               Tsf1SPILL10_256 <= Tspr10_2_V_1;
                               end 
                               end 
                      endcase
              if (!(!Tsf0SPILL14_256)) 
                  case (xpc10)
                      10'sd261/*261:xpc10*/:  begin 
                           xpc10 <= 10'sd195/*195:xpc10*/;
                           dfsin_gloops <= 32'sd1+dfsin_gloops;
                           end 
                          
                      10'sd263/*263:xpc10*/:  begin 
                           xpc10 <= 10'sd195/*195:xpc10*/;
                           dfsin_gloops <= 32'sd1+dfsin_gloops;
                           end 
                          endcase
                   else 
                  case (xpc10)
                      10'sd261/*261:xpc10*/:  begin 
                           xpc10 <= 10'sd247/*247:xpc10*/;
                           Tdbm0_3_V_2 <= Tdsi3_5_V_0;
                           end 
                          
                      10'sd263/*263:xpc10*/:  begin 
                           xpc10 <= 10'sd247/*247:xpc10*/;
                           Tdbm0_3_V_2 <= Tdsi3_5_V_0;
                           end 
                          endcase

              case (xpc10)
                  10'sd192/*192:xpc10*/:  begin 
                      if (!Tspr4_3_V_2 && !Tspr4_3_V_4 && !Tspr4_3_V_3)  begin 
                               xpc10 <= 10'sd193/*193:xpc10*/;
                               Tsf0_SPILL_256 <= Tspr4_3_V_0;
                               end 
                              if (!Tspr4_3_V_2 && !Tspr4_3_V_4 && Tspr4_3_V_3)  begin 
                               xpc10 <= 10'sd193/*193:xpc10*/;
                               Tsf0_SPILL_256 <= Tspr4_3_V_1;
                               end 
                              if (Tspr4_3_V_2 && !Tspr4_3_V_4)  begin 
                               xpc10 <= 10'sd193/*193:xpc10*/;
                               Tsf0_SPILL_256 <= Tspr4_3_V_0;
                               end 
                              if (Tspr4_3_V_4)  begin 
                               xpc10 <= 10'sd193/*193:xpc10*/;
                               Tsf0_SPILL_256 <= Tspr4_3_V_1;
                               end 
                               end 
                      
                  10'sd210/*210:xpc10*/:  begin 
                      if (!Tspr4_3_V_2 && !Tspr4_3_V_4 && !Tspr4_3_V_3)  begin 
                               xpc10 <= 10'sd211/*211:xpc10*/;
                               Tsf1_SPILL_256 <= Tspr4_3_V_0;
                               end 
                              if (!Tspr4_3_V_2 && !Tspr4_3_V_4 && Tspr4_3_V_3)  begin 
                               xpc10 <= 10'sd211/*211:xpc10*/;
                               Tsf1_SPILL_256 <= Tspr4_3_V_1;
                               end 
                              if (Tspr4_3_V_2 && !Tspr4_3_V_4)  begin 
                               xpc10 <= 10'sd211/*211:xpc10*/;
                               Tsf1_SPILL_256 <= Tspr4_3_V_0;
                               end 
                              if (Tspr4_3_V_4)  begin 
                               xpc10 <= 10'sd211/*211:xpc10*/;
                               Tsf1_SPILL_256 <= Tspr4_3_V_1;
                               end 
                               end 
                      
                  10'sd225/*225:xpc10*/:  begin 
                      if (!Tspr2_2_V_2 && !Tspr2_2_V_4 && !Tspr2_2_V_3)  begin 
                               xpc10 <= 10'sd226/*226:xpc10*/;
                               Tsf1SPILL10_256 <= Tspr2_2_V_0;
                               end 
                              if (!Tspr2_2_V_2 && !Tspr2_2_V_4 && Tspr2_2_V_3)  begin 
                               xpc10 <= 10'sd226/*226:xpc10*/;
                               Tsf1SPILL10_256 <= Tspr2_2_V_1;
                               end 
                              if (Tspr2_2_V_2 && !Tspr2_2_V_4)  begin 
                               xpc10 <= 10'sd226/*226:xpc10*/;
                               Tsf1SPILL10_256 <= Tspr2_2_V_0;
                               end 
                              if (Tspr2_2_V_4)  begin 
                               xpc10 <= 10'sd226/*226:xpc10*/;
                               Tsf1SPILL10_256 <= Tspr2_2_V_1;
                               end 
                               end 
                      
                  10'sd242/*242:xpc10*/:  begin 
                      if (!Tspr3_2_V_2 && !Tspr3_2_V_4 && !Tspr3_2_V_3)  begin 
                               xpc10 <= 10'sd243/*243:xpc10*/;
                               Tsa1_SPILL_256 <= Tspr3_2_V_0;
                               end 
                              if (!Tspr3_2_V_2 && !Tspr3_2_V_4 && Tspr3_2_V_3)  begin 
                               xpc10 <= 10'sd243/*243:xpc10*/;
                               Tsa1_SPILL_256 <= Tspr3_2_V_1;
                               end 
                              if (Tspr3_2_V_2 && !Tspr3_2_V_4)  begin 
                               xpc10 <= 10'sd243/*243:xpc10*/;
                               Tsa1_SPILL_256 <= Tspr3_2_V_0;
                               end 
                              if (Tspr3_2_V_4)  begin 
                               xpc10 <= 10'sd243/*243:xpc10*/;
                               Tsa1_SPILL_256 <= Tspr3_2_V_1;
                               end 
                               end 
                      endcase
              if (!Tspr4_3_V_2 && !Tspr4_3_V_4 && !Tspr4_3_V_3) 
                  case (xpc10)
                      10'sd191/*191:xpc10*/:  begin 
                           xpc10 <= 10'sd193/*193:xpc10*/;
                           Tsf0_SPILL_256 <= Tspr4_3_V_0;
                           end 
                          
                      10'sd209/*209:xpc10*/:  begin 
                           xpc10 <= 10'sd211/*211:xpc10*/;
                           Tsf1_SPILL_256 <= Tspr4_3_V_0;
                           end 
                          endcase
                  if (!Tspr4_3_V_2 && !Tspr4_3_V_4 && Tspr4_3_V_3) 
                  case (xpc10)
                      10'sd191/*191:xpc10*/:  begin 
                           xpc10 <= 10'sd193/*193:xpc10*/;
                           Tsf0_SPILL_256 <= Tspr4_3_V_1;
                           end 
                          
                      10'sd209/*209:xpc10*/:  begin 
                           xpc10 <= 10'sd211/*211:xpc10*/;
                           Tsf1_SPILL_256 <= Tspr4_3_V_1;
                           end 
                          endcase
                  if ((64'sh0<(A_64_US_CC_SCALbx12_ARB0[Tdbm0_3_V_1]>>32'sd63))) 
                  case (xpc10)
                      10'sd179/*179:xpc10*/:  begin 
                           xpc10 <= 10'sd180/*180:xpc10*/;
                           Tsfl0_9_V_0 <= 1'h1;
                           end 
                          
                      10'sd182/*182:xpc10*/:  begin 
                           xpc10 <= 10'sd183/*183:xpc10*/;
                           Tsfl0_9_V_1 <= 1'h1;
                           end 
                          endcase
                   else 
                  case (xpc10)
                      10'sd179/*179:xpc10*/:  begin 
                           xpc10 <= 10'sd180/*180:xpc10*/;
                           Tsfl0_9_V_0 <= 1'h0;
                           end 
                          
                      10'sd182/*182:xpc10*/:  begin 
                           xpc10 <= 10'sd183/*183:xpc10*/;
                           Tsfl0_9_V_1 <= 1'h0;
                           end 
                          endcase
              if ((xpc10==10'sd253/*253:xpc10*/))  begin 
                      if ((Tdbm0_3_V_0!=32'sd36/*36:Tdbm0.3_V_0*/) && (Tdbm0_3_V_1>=32'sd36))  xpc10 <= 10'sd256/*256:xpc10*/;
                          if ((Tdbm0_3_V_0==32'sd36/*36:Tdbm0.3_V_0*/) && (Tdbm0_3_V_1>=32'sd36))  xpc10 <= 10'sd254/*254:xpc10*/;
                          if ((Tdbm0_3_V_1<32'sd36))  xpc10 <= 10'sd174/*174:xpc10*/;
                           end 
                      if ((Tsfl0_9_V_9==32'sd0/*0:Tsfl0.9_V_9*/))  begin if ((xpc10==10'sd790/*790:xpc10*/))  begin 
                           xpc10 <= 10'sd822/*822:xpc10*/;
                           Tsf0_SPILL_259 <= 64'sh0;
                           Tsf0_SPILL_257 <= fastspilldup20;
                           end 
                           end 
                   else if ((xpc10==10'sd790/*790:xpc10*/))  begin 
                           xpc10 <= 10'sd791/*791:xpc10*/;
                           Tsf0_SPILL_259 <= 64'sh1;
                           Tsf0_SPILL_257 <= fastspilldup20;
                           end 
                          if ((Tsfl1_7_V_9==32'sd0/*0:Tsfl1.7_V_9*/))  begin if ((xpc10==10'sd692/*692:xpc10*/))  begin 
                           xpc10 <= 10'sd724/*724:xpc10*/;
                           Tsf1_SPILL_259 <= 64'sh0;
                           Tsf1_SPILL_257 <= fastspilldup30;
                           end 
                           end 
                   else if ((xpc10==10'sd692/*692:xpc10*/))  begin 
                           xpc10 <= 10'sd693/*693:xpc10*/;
                           Tsf1_SPILL_259 <= 64'sh1;
                           Tsf1_SPILL_257 <= fastspilldup30;
                           end 
                          
              case (xpc10)
                  10'sd567/*567:xpc10*/: if ((Tsad27_13_V_0<Tsfl1_18_V_10))  begin 
                           xpc10 <= 10'sd568/*568:xpc10*/;
                           Tsa27_SPILL_259 <= Tsa27_SPILL_257;
                           Tsa27_SPILL_260 <= 64'sh1;
                           end 
                           else  begin 
                           xpc10 <= 10'sd570/*570:xpc10*/;
                           Tsa27_SPILL_259 <= Tsa27_SPILL_262;
                           Tsa27_SPILL_260 <= 64'sh0;
                           end 
                          
                  10'sd586/*586:xpc10*/: if ((Tsmu5_7_V_5<Tsmu5_7_V_6))  begin 
                           xpc10 <= 10'sd587/*587:xpc10*/;
                           Tsm5_SPILL_259 <= 64'sh1;
                           Tsm5_SPILL_257 <= fastspilldup36;
                           end 
                           else  begin 
                           xpc10 <= 10'sd615/*615:xpc10*/;
                           Tsm5_SPILL_259 <= 64'sh0;
                           Tsm5_SPILL_257 <= fastspilldup36;
                           end 
                          
                  10'sd591/*591:xpc10*/: if ((Tsmu5_7_V_7<Tsmu5_7_V_5))  begin 
                           xpc10 <= 10'sd592/*592:xpc10*/;
                           Tsm5_SPILL_262 <= 64'sh1;
                           Tsm5_SPILL_260 <= fastspilldup38;
                           end 
                           else  begin 
                           xpc10 <= 10'sd614/*614:xpc10*/;
                           Tsm5_SPILL_262 <= 64'sh0;
                           Tsm5_SPILL_260 <= fastspilldup38;
                           end 
                          
                  10'sd597/*597:xpc10*/: if ((64'sh0<Tses25_5_V_5))  begin 
                           xpc10 <= 10'sd598/*598:xpc10*/;
                           Tss5_SPILL_259 <= Tss5_SPILL_257;
                           Tss5_SPILL_260 <= 64'sh1;
                           end 
                           else  begin 
                           xpc10 <= 10'sd613/*613:xpc10*/;
                           Tss5_SPILL_259 <= Tss5_SPILL_262;
                           Tss5_SPILL_260 <= 64'sh0;
                           end 
                          
                  10'sd601/*601:xpc10*/: if ((Tses25_5_V_2<(Tses25_5_V_0<<32'sd32)))  begin 
                           xpc10 <= 10'sd604/*604:xpc10*/;
                           Tse25_SPILL_260 <= (Tses25_5_V_2/Tses25_5_V_0);
                           Tse25_SPILL_258 <= fastspilldup44;
                           end 
                           else  begin 
                           xpc10 <= 10'sd602/*602:xpc10*/;
                           Tse25_SPILL_260 <= 64'h_ffff_ffff;
                           Tse25_SPILL_258 <= fastspilldup44;
                           end 
                          
                  10'sd609/*609:xpc10*/: if ((Tsad6_15_V_0<Tses25_5_V_3))  begin 
                           xpc10 <= 10'sd610/*610:xpc10*/;
                           Tsa6_SPILL_259 <= Tsa6_SPILL_257;
                           Tsa6_SPILL_260 <= 64'sh1;
                           end 
                           else  begin 
                           xpc10 <= 10'sd612/*612:xpc10*/;
                           Tsa6_SPILL_259 <= Tsa6_SPILL_262;
                           Tsa6_SPILL_260 <= 64'sh0;
                           end 
                          endcase
              if ((32'sd0/*0:USA74*/==(Tsro33_4_V_1<<(32'sd63&rtl_signed_bitextract0(Tsro33_4_V_0)))))  begin if ((xpc10==10'sd556/*556:xpc10*/)) 
                   begin 
                           xpc10 <= 10'sd559/*559:xpc10*/;
                           Tss18_SPILL_257 <= Tss18_SPILL_259;
                           Tss18_SPILL_258 <= 64'sh0;
                           end 
                           end 
                   else if ((xpc10==10'sd556/*556:xpc10*/))  begin 
                           xpc10 <= 10'sd557/*557:xpc10*/;
                           Tss18_SPILL_257 <= Tss18_SPILL_256;
                           Tss18_SPILL_258 <= 64'sh1;
                           end 
                          if (!(!Tsro33_4_V_6)) 
                  case (xpc10)
                      10'sd547/*547:xpc10*/:  xpc10 <= 10'sd548/*548:xpc10*/;

                      10'sd548/*548:xpc10*/:  xpc10 <= 10'sd549/*549:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      10'sd547/*547:xpc10*/:  begin 
                           xpc10 <= 10'sd550/*550:xpc10*/;
                           Tsro33_4_V_1 <= (Tsro33_4_V_1+rtl_sign_extend4(Tsro33_4_V_5)>>32'sd10);
                           end 
                          
                      10'sd548/*548:xpc10*/:  begin 
                           xpc10 <= 10'sd550/*550:xpc10*/;
                           Tsro33_4_V_1 <= (Tsro33_4_V_1+rtl_sign_extend4(Tsro33_4_V_5)>>32'sd10);
                           end 
                          endcase
              if ((xpc10==10'sd541/*541:xpc10*/)) if (!(!Tsro33_4_V_5))  begin 
                           xpc10 <= 10'sd544/*544:xpc10*/;
                           Tsr33_SPILL_257 <= Tsr33_SPILL_260;
                           Tsr33_SPILL_258 <= 64'sh0;
                           end 
                           else  begin 
                           xpc10 <= 10'sd542/*542:xpc10*/;
                           Tsr33_SPILL_257 <= Tsr33_SPILL_256;
                           Tsr33_SPILL_258 <= 64'sh1;
                           end 
                          if ((Tsfl1_18_V_10==32'sd0/*0:Tsfl1.18_V_10*/))  begin if ((xpc10==10'sd533/*533:xpc10*/))  begin 
                           xpc10 <= 10'sd563/*563:xpc10*/;
                           Tsf1SPILL10_259 <= 64'sh0;
                           Tsf1SPILL10_257 <= fastspilldup54;
                           end 
                           end 
                   else if ((xpc10==10'sd533/*533:xpc10*/))  begin 
                           xpc10 <= 10'sd534/*534:xpc10*/;
                           Tsf1SPILL10_259 <= 64'sh1;
                           Tsf1SPILL10_257 <= fastspilldup54;
                           end 
                          
              case (xpc10)
                  10'sd447/*447:xpc10*/:  begin 
                      if ((Tssu2_4_V_5>=Tssu2_4_V_4) && (Tssu2_4_V_4>=Tssu2_4_V_5))  begin 
                               xpc10 <= 10'sd448/*448:xpc10*/;
                               Tss2_SPILL_256 <= 64'h0;
                               end 
                              if ((Tssu2_4_V_5>=Tssu2_4_V_4) && (Tssu2_4_V_4<Tssu2_4_V_5))  begin 
                               xpc10 <= 10'sd427/*427:xpc10*/;
                               Tssu2_4_V_6 <= Tssu2_4_V_5+(0-Tssu2_4_V_4);
                               end 
                              if ((Tssu2_4_V_5<Tssu2_4_V_4))  begin 
                               xpc10 <= 10'sd367/*367:xpc10*/;
                               Tssu2_4_V_6 <= Tssu2_4_V_4+(0-Tssu2_4_V_5);
                               end 
                               end 
                      
                  10'sd449/*449:xpc10*/:  begin 
                      if ((Tsfl1_22_V_0? !rtl_unsigned_bitextract5(Tse0SPILL18_256): rtl_unsigned_bitextract5(Tse0SPILL18_256)))  begin 
                               xpc10 <= 10'sd345/*345:xpc10*/;
                               Tssu2_4_V_0 <= rtl_unsigned_bitextract8(Tsfl1_22_V_0);
                               Tsfl1_22_V_1 <= rtl_unsigned_bitextract5(Tse0SPILL18_256);
                               end 
                              if ((Tsfl1_22_V_0? rtl_unsigned_bitextract5(Tse0SPILL18_256): !rtl_unsigned_bitextract5(Tse0SPILL18_256
                      )))  begin 
                               xpc10 <= 10'sd229/*229:xpc10*/;
                               Tsad1_3_V_3 <= 64'shf_ffff_ffff_ffff&Tdsi3_5_V_0;
                               Tsfl1_22_V_1 <= rtl_unsigned_bitextract5(Tse0SPILL18_256);
                               end 
                               end 
                      
                  10'sd505/*505:xpc10*/:  begin 
                      if ((Tsfl1_18_V_6+Tsfl1_18_V_6<Tsfl1_18_V_7) && (Tsfl1_18_V_6<Tsfl1_18_V_7))  begin 
                               xpc10 <= 10'sd574/*574:xpc10*/;
                               Tses25_5_V_0 <= (Tsfl1_18_V_7>>32'sd32);
                               end 
                              if ((Tsfl1_18_V_6+Tsfl1_18_V_6<Tsfl1_18_V_7) && (Tsfl1_18_V_6>=Tsfl1_18_V_7))  begin 
                               xpc10 <= 10'sd508/*508:xpc10*/;
                               Tsfl1_18_V_8 <= 64'h_ffff_ffff_ffff_ffff;
                               end 
                              if ((Tsfl1_18_V_6+Tsfl1_18_V_6>=Tsfl1_18_V_7))  begin 
                               xpc10 <= 10'sd506/*506:xpc10*/;
                               Tsfl1_18_V_6 <= (Tsfl1_18_V_6>>32'sd1);
                               end 
                               end 
                      
                  10'sd519/*519:xpc10*/: if ((Tsmu26_4_V_5<Tsmu26_4_V_6))  begin 
                           xpc10 <= 10'sd520/*520:xpc10*/;
                           Tsm26_SPILL_259 <= 64'sh1;
                           Tsm26_SPILL_257 <= fastspilldup46;
                           end 
                           else  begin 
                           xpc10 <= 10'sd573/*573:xpc10*/;
                           Tsm26_SPILL_259 <= 64'sh0;
                           Tsm26_SPILL_257 <= fastspilldup46;
                           end 
                          
                  10'sd524/*524:xpc10*/: if ((Tsmu26_4_V_7<Tsmu26_4_V_5))  begin 
                           xpc10 <= 10'sd525/*525:xpc10*/;
                           Tsm26_SPILL_262 <= 64'sh1;
                           Tsm26_SPILL_260 <= fastspilldup48;
                           end 
                           else  begin 
                           xpc10 <= 10'sd572/*572:xpc10*/;
                           Tsm26_SPILL_262 <= 64'sh0;
                           Tsm26_SPILL_260 <= fastspilldup48;
                           end 
                          
                  10'sd530/*530:xpc10*/: if ((64'sh0<Tsfl1_18_V_12))  begin 
                           xpc10 <= 10'sd531/*531:xpc10*/;
                           Tss26_SPILL_259 <= Tss26_SPILL_257;
                           Tss26_SPILL_260 <= 64'sh1;
                           end 
                           else  begin 
                           xpc10 <= 10'sd571/*571:xpc10*/;
                           Tss26_SPILL_259 <= Tss26_SPILL_262;
                           Tss26_SPILL_260 <= 64'sh0;
                           end 
                          endcase
              if ((32'sd0/*0:USA148*/==(Tssu2_4_V_4<<(32'sd63&rtl_signed_bitextract0(Tssu2_4_V_7)))))  begin if ((xpc10==10'sd430/*430:xpc10*/)) 
                   begin 
                           xpc10 <= 10'sd433/*433:xpc10*/;
                           Tss23_SPILL_257 <= Tss23_SPILL_259;
                           Tss23_SPILL_258 <= 64'sh0;
                           end 
                           end 
                   else if ((xpc10==10'sd430/*430:xpc10*/))  begin 
                           xpc10 <= 10'sd431/*431:xpc10*/;
                           Tss23_SPILL_257 <= Tss23_SPILL_256;
                           Tss23_SPILL_258 <= 64'sh1;
                           end 
                          if ((32'sd0/*0:USA134*/==(Tssu2_4_V_5<<(32'sd63&rtl_signed_bitextract0((0-Tssu2_4_V_7))))))  begin if ((xpc10
                  ==10'sd407/*407:xpc10*/))  begin 
                           xpc10 <= 10'sd410/*410:xpc10*/;
                           Tss32_SPILL_257 <= Tss32_SPILL_259;
                           Tss32_SPILL_258 <= 64'sh0;
                           end 
                           end 
                   else if ((xpc10==10'sd407/*407:xpc10*/))  begin 
                           xpc10 <= 10'sd408/*408:xpc10*/;
                           Tss32_SPILL_257 <= Tss32_SPILL_256;
                           Tss32_SPILL_258 <= 64'sh1;
                           end 
                          if ((32'sd0/*0:USA162*/==(Tsro0_16_V_1<<(32'sd63&rtl_signed_bitextract0(Tsro0_16_V_0)))))  begin if ((xpc10
                  ==10'sd398/*398:xpc10*/))  begin 
                           xpc10 <= 10'sd401/*401:xpc10*/;
                           Tss18_SPILL_257 <= Tss18_SPILL_259;
                           Tss18_SPILL_258 <= 64'sh0;
                           end 
                           end 
                   else if ((xpc10==10'sd398/*398:xpc10*/))  begin 
                           xpc10 <= 10'sd399/*399:xpc10*/;
                           Tss18_SPILL_257 <= Tss18_SPILL_256;
                           Tss18_SPILL_258 <= 64'sh1;
                           end 
                          if (!(!Tsro0_16_V_6)) 
                  case (xpc10)
                      10'sd389/*389:xpc10*/:  xpc10 <= 10'sd390/*390:xpc10*/;

                      10'sd390/*390:xpc10*/:  xpc10 <= 10'sd391/*391:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      10'sd389/*389:xpc10*/:  begin 
                           xpc10 <= 10'sd392/*392:xpc10*/;
                           Tsro0_16_V_1 <= (Tsro0_16_V_1+rtl_sign_extend4(Tsro0_16_V_5)>>32'sd10);
                           end 
                          
                      10'sd390/*390:xpc10*/:  begin 
                           xpc10 <= 10'sd392/*392:xpc10*/;
                           Tsro0_16_V_1 <= (Tsro0_16_V_1+rtl_sign_extend4(Tsro0_16_V_5)>>32'sd10);
                           end 
                          endcase
              if ((xpc10==10'sd383/*383:xpc10*/)) if (!(!Tsro0_16_V_5))  begin 
                           xpc10 <= 10'sd386/*386:xpc10*/;
                           Tsr0_SPILL_257 <= Tsr0_SPILL_260;
                           Tsr0_SPILL_258 <= 64'sh0;
                           end 
                           else  begin 
                           xpc10 <= 10'sd384/*384:xpc10*/;
                           Tsr0_SPILL_257 <= Tsr0_SPILL_256;
                           Tsr0_SPILL_258 <= 64'sh1;
                           end 
                          if ((32'sd0/*0:USA104*/==(Tsad1_3_V_3<<(32'sd63&rtl_signed_bitextract0(Tsad1_3_V_6)))))  begin if ((xpc10==
                  10'sd323/*323:xpc10*/))  begin 
                           xpc10 <= 10'sd327/*327:xpc10*/;
                           Tss17_SPILL_257 <= Tss17_SPILL_259;
                           Tss17_SPILL_258 <= 64'sh0;
                           end 
                           end 
                   else if ((xpc10==10'sd323/*323:xpc10*/))  begin 
                           xpc10 <= 10'sd324/*324:xpc10*/;
                           Tss17_SPILL_257 <= Tss17_SPILL_256;
                           Tss17_SPILL_258 <= 64'sh1;
                           end 
                          if ((32'sd0/*0:USA90*/==(Tsad1_3_V_4<<(32'sd63&rtl_signed_bitextract0((0-Tsad1_3_V_6))))))  begin if ((xpc10
                  ==10'sd302/*302:xpc10*/))  begin 
                           xpc10 <= 10'sd306/*306:xpc10*/;
                           Tss8_SPILL_257 <= Tss8_SPILL_259;
                           Tss8_SPILL_258 <= 64'sh0;
                           end 
                           end 
                   else if ((xpc10==10'sd302/*302:xpc10*/))  begin 
                           xpc10 <= 10'sd303/*303:xpc10*/;
                           Tss8_SPILL_257 <= Tss8_SPILL_256;
                           Tss8_SPILL_258 <= 64'sh1;
                           end 
                          if ((32'sd0/*0:USA118*/==(Tsro28_4_V_1<<(32'sd63&rtl_signed_bitextract0(Tsro28_4_V_0)))))  begin if ((xpc10
                  ==10'sd294/*294:xpc10*/))  begin 
                           xpc10 <= 10'sd297/*297:xpc10*/;
                           Tss18_SPILL_257 <= Tss18_SPILL_259;
                           Tss18_SPILL_258 <= 64'sh0;
                           end 
                           end 
                   else if ((xpc10==10'sd294/*294:xpc10*/))  begin 
                           xpc10 <= 10'sd295/*295:xpc10*/;
                           Tss18_SPILL_257 <= Tss18_SPILL_256;
                           Tss18_SPILL_258 <= 64'sh1;
                           end 
                          if (!(!Tsro28_4_V_6)) 
                  case (xpc10)
                      10'sd285/*285:xpc10*/:  xpc10 <= 10'sd286/*286:xpc10*/;

                      10'sd286/*286:xpc10*/:  xpc10 <= 10'sd287/*287:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      10'sd285/*285:xpc10*/:  begin 
                           xpc10 <= 10'sd288/*288:xpc10*/;
                           Tsro28_4_V_1 <= (Tsro28_4_V_1+rtl_sign_extend4(Tsro28_4_V_5)>>32'sd10);
                           end 
                          
                      10'sd286/*286:xpc10*/:  begin 
                           xpc10 <= 10'sd288/*288:xpc10*/;
                           Tsro28_4_V_1 <= (Tsro28_4_V_1+rtl_sign_extend4(Tsro28_4_V_5)>>32'sd10);
                           end 
                          endcase

              case (xpc10)
                  10'sd260/*260:xpc10*/: if (!(!Tsf0SPILL14_257))  begin 
                           xpc10 <= 10'sd195/*195:xpc10*/;
                           dfsin_gloops <= 32'sd1+dfsin_gloops;
                           Tsf0SPILL14_256 <= Tsf0SPILL14_257;
                           end 
                           else  begin 
                           xpc10 <= 10'sd247/*247:xpc10*/;
                           Tdbm0_3_V_2 <= Tdsi3_5_V_0;
                           Tsf0SPILL14_256 <= Tsf0SPILL14_257;
                           end 
                          
                  10'sd262/*262:xpc10*/: if (!(!Tsf0SPILL14_258))  begin 
                           xpc10 <= 10'sd195/*195:xpc10*/;
                           dfsin_gloops <= 32'sd1+dfsin_gloops;
                           Tsf0SPILL14_256 <= Tsf0SPILL14_258;
                           end 
                           else  begin 
                           xpc10 <= 10'sd247/*247:xpc10*/;
                           Tdbm0_3_V_2 <= Tdsi3_5_V_0;
                           Tsf0SPILL14_256 <= Tsf0SPILL14_258;
                           end 
                          
                  10'sd279/*279:xpc10*/: if (!(!Tsro28_4_V_5))  begin 
                           xpc10 <= 10'sd282/*282:xpc10*/;
                           Tsr28_SPILL_257 <= Tsr28_SPILL_260;
                           Tsr28_SPILL_258 <= 64'sh0;
                           end 
                           else  begin 
                           xpc10 <= 10'sd280/*280:xpc10*/;
                           Tsr28_SPILL_257 <= Tsr28_SPILL_256;
                           Tsr28_SPILL_258 <= 64'sh1;
                           end 
                          endcase
              if ((Tdbm0_3_V_2==A_64_US_CC_SCALbx10_ARA0[Tdbm0_3_V_1]))  begin if ((xpc10==10'sd248/*248:xpc10*/))  begin 
                           xpc10 <= 10'sd249/*249:xpc10*/;
                           Tdb0_SPILL_258 <= 32'sd1;
                           Tdb0_SPILL_256 <= fastspilldup76;
                           end 
                           end 
                   else if ((xpc10==10'sd248/*248:xpc10*/))  begin 
                           xpc10 <= 10'sd257/*257:xpc10*/;
                           Tdb0_SPILL_258 <= 32'sd0;
                           Tdb0_SPILL_256 <= fastspilldup76;
                           end 
                          if ((Tsfl1_22_V_0? (xpc10==10'sd228/*228:xpc10*/) && !rtl_unsigned_bitextract5(Tse0SPILL18_256): (xpc10==10'sd228
              /*228:xpc10*/) && rtl_unsigned_bitextract5(Tse0SPILL18_256)))  begin 
                       xpc10 <= 10'sd345/*345:xpc10*/;
                       Tssu2_4_V_0 <= rtl_unsigned_bitextract8(Tsfl1_22_V_0);
                       Tsfl1_22_V_1 <= rtl_unsigned_bitextract5(Tse0SPILL18_256);
                       end 
                      if ((Tsfl1_22_V_0? (xpc10==10'sd228/*228:xpc10*/) && rtl_unsigned_bitextract5(Tse0SPILL18_256): (xpc10==10'sd228
              /*228:xpc10*/) && !rtl_unsigned_bitextract5(Tse0SPILL18_256)))  begin 
                       xpc10 <= 10'sd229/*229:xpc10*/;
                       Tsad1_3_V_3 <= 64'shf_ffff_ffff_ffff&Tdsi3_5_V_0;
                       Tsfl1_22_V_1 <= rtl_unsigned_bitextract5(Tse0SPILL18_256);
                       end 
                      if ((xpc10==10'sd792/*792:xpc10*/)) if (($signed((Tsfl0_9_V_8<<32'sd1))<64'sh0))  begin 
                           xpc10 <= 10'sd795/*795:xpc10*/;
                           Tsro29_4_V_1 <= Tsfl0_9_V_8;
                           Tsro29_4_V_0 <= rtl_signed_bitextract0(Tsfl0_9_V_5);
                           end 
                           else  begin 
                           xpc10 <= 10'sd793/*793:xpc10*/;
                           Tsfl0_9_V_8 <= (Tsfl0_9_V_8<<32'sd1);
                           end 
                          if ((Tspr11_2_V_2 || Tspr11_2_V_4) && (xpc10==10'sd739/*739:xpc10*/))  xpc10 <= 10'sd740/*740:xpc10*/;
                  if ((xpc10==10'sd694/*694:xpc10*/)) if (($signed((Tsfl1_7_V_8<<32'sd1))<64'sh0))  begin 
                           xpc10 <= 10'sd697/*697:xpc10*/;
                           Tsro29_4_V_1 <= Tsfl1_7_V_8;
                           Tsro29_4_V_0 <= rtl_signed_bitextract0(Tsfl1_7_V_5);
                           end 
                           else  begin 
                           xpc10 <= 10'sd695/*695:xpc10*/;
                           Tsfl1_7_V_8 <= (Tsfl1_7_V_8<<32'sd1);
                           end 
                          if ((Tspr11_2_V_2 || Tspr11_2_V_4) && (xpc10==10'sd641/*641:xpc10*/))  xpc10 <= 10'sd642/*642:xpc10*/;
                  
              case (xpc10)
                  10'sd473/*473:xpc10*/:  begin 
                      if (!Tspr10_2_V_2 && !Tspr10_2_V_4 && !Tspr10_2_V_3)  begin 
                               xpc10 <= 10'sd475/*475:xpc10*/;
                               Tsf1SPILL10_256 <= Tspr10_2_V_0;
                               end 
                              if (!Tspr10_2_V_2 && !Tspr10_2_V_4 && Tspr10_2_V_3)  begin 
                               xpc10 <= 10'sd475/*475:xpc10*/;
                               Tsf1SPILL10_256 <= Tspr10_2_V_1;
                               end 
                              if (Tspr10_2_V_2 || Tspr10_2_V_4)  begin if (Tspr10_2_V_2 || Tspr10_2_V_4)  xpc10 <= 10'sd474/*474:xpc10*/;
                               end 
                           end 
                      
                  10'sd508/*508:xpc10*/: if ((64'sh2<(64'sh1ff&Tsfl1_18_V_8)))  begin 
                           xpc10 <= 10'sd536/*536:xpc10*/;
                           Tsro33_4_V_1 <= Tsfl1_18_V_8;
                           Tsro33_4_V_0 <= rtl_signed_bitextract0(Tsfl1_18_V_5);
                           end 
                           else  begin 
                           xpc10 <= 10'sd509/*509:xpc10*/;
                           Tsmu26_4_V_1 <= rtl_unsigned_bitextract1(64'h_ffff_ffff&Tsfl1_18_V_7);
                           end 
                          
                  10'sd574/*574:xpc10*/: if ((Tsfl1_18_V_6<(Tses25_5_V_0<<32'sd32)))  begin 
                           xpc10 <= 10'sd616/*616:xpc10*/;
                           Tse25_SPILL_257 <= ((Tsfl1_18_V_6/Tses25_5_V_0)<<32'sd32);
                           end 
                           else  begin 
                           xpc10 <= 10'sd575/*575:xpc10*/;
                           Tses25_5_V_6 <= 64'h_ffff_ffff_0000_0000;
                           Tse25_SPILL_257 <= 64'h_ffff_ffff_0000_0000;
                           end 
                          endcase
              if ((32'sd4094/*4094:USA68*/==(64'shfff&(Tspr10_2_V_1>>32'sd51))))  begin if ((xpc10==10'sd470/*470:xpc10*/))  begin 
                           xpc10 <= 10'sd471/*471:xpc10*/;
                           Tsf0SPILL12_256 <= rtl_sign_extend6((32'sd0/*0:USA72*/==(32'sd0/*0:USA70*/==(64'sh7_ffff_ffff_ffff&Tspr10_2_V_1
                          ))));

                           end 
                           end 
                   else if ((xpc10==10'sd470/*470:xpc10*/))  begin 
                           xpc10 <= 10'sd476/*476:xpc10*/;
                           Tspr10_2_V_4 <= 1'h0;
                           Tsf0SPILL12_256 <= 32'sd0;
                           end 
                          if ((32'sd4094/*4094:USA62*/==(64'shfff&(Tspr10_2_V_0>>32'sd51))))  begin if ((xpc10==10'sd468/*468:xpc10*/)) 
                   begin 
                           xpc10 <= 10'sd469/*469:xpc10*/;
                           Tsf0SPILL10_256 <= rtl_sign_extend6((32'sd0/*0:USA66*/==(32'sd0/*0:USA64*/==(64'sh7_ffff_ffff_ffff&Tspr10_2_V_0
                          ))));

                           end 
                           end 
                   else if ((xpc10==10'sd468/*468:xpc10*/))  begin 
                           xpc10 <= 10'sd477/*477:xpc10*/;
                           Tspr10_2_V_2 <= 1'h0;
                           Tsf0SPILL10_256 <= 32'sd0;
                           end 
                          
              case (xpc10)
                  10'sd458/*458:xpc10*/:  begin 
                      if (!Tspr5_2_V_2 && !Tspr5_2_V_4 && !Tspr5_2_V_3)  begin 
                               xpc10 <= 10'sd460/*460:xpc10*/;
                               Tsf1SPILL10_256 <= Tspr5_2_V_0;
                               end 
                              if (!Tspr5_2_V_2 && !Tspr5_2_V_4 && Tspr5_2_V_3)  begin 
                               xpc10 <= 10'sd460/*460:xpc10*/;
                               Tsf1SPILL10_256 <= Tspr5_2_V_1;
                               end 
                              if (Tspr5_2_V_2 || Tspr5_2_V_4)  begin if (Tspr5_2_V_2 || Tspr5_2_V_4)  xpc10 <= 10'sd459/*459:xpc10*/;
                               end 
                           end 
                      
                  10'sd466/*466:xpc10*/:  begin 
                      if ((Tsfl1_22_V_0? !Tsfl1_22_V_1: Tsfl1_22_V_1))  begin 
                               xpc10 <= 10'sd346/*346:xpc10*/;
                               Tssu2_4_V_4 <= 64'shf_ffff_ffff_ffff&Tdsi3_5_V_0;
                               Tssu2_4_V_0 <= rtl_unsigned_bitextract8(Tsfl1_22_V_0);
                               end 
                              if ((Tsfl1_22_V_0? Tsfl1_22_V_1: !Tsfl1_22_V_1))  begin 
                               xpc10 <= 10'sd229/*229:xpc10*/;
                               Tsad1_3_V_3 <= 64'shf_ffff_ffff_ffff&Tdsi3_5_V_0;
                               end 
                               end 
                      endcase
              if ((32'sd4094/*4094:USA56*/==(64'shfff&(Tspr5_2_V_1>>32'sd51))))  begin if ((xpc10==10'sd455/*455:xpc10*/))  begin 
                           xpc10 <= 10'sd456/*456:xpc10*/;
                           Tsf0SPILL12_256 <= rtl_sign_extend6((32'sd0/*0:USA60*/==(32'sd0/*0:USA58*/==(64'sh7_ffff_ffff_ffff&Tspr5_2_V_1
                          ))));

                           end 
                           end 
                   else if ((xpc10==10'sd455/*455:xpc10*/))  begin 
                           xpc10 <= 10'sd461/*461:xpc10*/;
                           Tspr5_2_V_4 <= 1'h0;
                           Tsf0SPILL12_256 <= 32'sd0;
                           end 
                          if ((32'sd4094/*4094:USA50*/==(64'shfff&(Tspr5_2_V_0>>32'sd51))))  begin if ((xpc10==10'sd453/*453:xpc10*/)) 
                   begin 
                           xpc10 <= 10'sd454/*454:xpc10*/;
                           Tsf0SPILL10_256 <= rtl_sign_extend6((32'sd0/*0:USA54*/==(32'sd0/*0:USA52*/==(64'sh7_ffff_ffff_ffff&Tspr5_2_V_0
                          ))));

                           end 
                           end 
                   else if ((xpc10==10'sd453/*453:xpc10*/))  begin 
                           xpc10 <= 10'sd462/*462:xpc10*/;
                           Tspr5_2_V_2 <= 1'h0;
                           Tsf0SPILL10_256 <= 32'sd0;
                           end 
                          if ((xpc10==10'sd441/*441:xpc10*/))  begin 
                      if (!Tspr7_3_V_2 && !Tspr7_3_V_4 && !Tspr7_3_V_3)  begin 
                               xpc10 <= 10'sd443/*443:xpc10*/;
                               Tss2_SPILL_256 <= Tspr7_3_V_0;
                               end 
                              if (!Tspr7_3_V_2 && !Tspr7_3_V_4 && Tspr7_3_V_3)  begin 
                               xpc10 <= 10'sd443/*443:xpc10*/;
                               Tss2_SPILL_256 <= Tspr7_3_V_1;
                               end 
                              if (Tspr7_3_V_2 || Tspr7_3_V_4)  begin if (Tspr7_3_V_2 || Tspr7_3_V_4)  xpc10 <= 10'sd442/*442:xpc10*/;
                               end 
                           end 
                      if ((32'sd4094/*4094:USA156*/==(64'shfff&(Tspr7_3_V_1>>32'sd51))))  begin if ((xpc10==10'sd438/*438:xpc10*/))  begin 
                           xpc10 <= 10'sd439/*439:xpc10*/;
                           Tsf0SPILL12_256 <= rtl_sign_extend6((32'sd0/*0:USA160*/==(32'sd0/*0:USA158*/==(64'sh7_ffff_ffff_ffff&Tspr7_3_V_1
                          ))));

                           end 
                           end 
                   else if ((xpc10==10'sd438/*438:xpc10*/))  begin 
                           xpc10 <= 10'sd444/*444:xpc10*/;
                           Tspr7_3_V_4 <= 1'h0;
                           Tsf0SPILL12_256 <= 32'sd0;
                           end 
                          if ((32'sd4094/*4094:USA150*/==(64'shfff&(Tspr7_3_V_0>>32'sd51))))  begin if ((xpc10==10'sd436/*436:xpc10*/)) 
                   begin 
                           xpc10 <= 10'sd437/*437:xpc10*/;
                           Tsf0SPILL10_256 <= rtl_sign_extend6((32'sd0/*0:USA154*/==(32'sd0/*0:USA152*/==(64'sh7_ffff_ffff_ffff&Tspr7_3_V_0
                          ))));

                           end 
                           end 
                   else if ((xpc10==10'sd436/*436:xpc10*/))  begin 
                           xpc10 <= 10'sd445/*445:xpc10*/;
                           Tspr7_3_V_2 <= 1'h0;
                           Tsf0SPILL10_256 <= 32'sd0;
                           end 
                          if ((xpc10==10'sd418/*418:xpc10*/))  begin 
                      if (!Tspr18_2_V_2 && !Tspr18_2_V_4 && !Tspr18_2_V_3)  begin 
                               xpc10 <= 10'sd420/*420:xpc10*/;
                               Tss2_SPILL_256 <= Tspr18_2_V_0;
                               end 
                              if (!Tspr18_2_V_2 && !Tspr18_2_V_4 && Tspr18_2_V_3)  begin 
                               xpc10 <= 10'sd420/*420:xpc10*/;
                               Tss2_SPILL_256 <= Tspr18_2_V_1;
                               end 
                              if (Tspr18_2_V_2 || Tspr18_2_V_4)  begin if (Tspr18_2_V_2 || Tspr18_2_V_4)  xpc10 <= 10'sd419/*419:xpc10*/;
                               end 
                           end 
                      if ((32'sd4094/*4094:USA142*/==(64'shfff&(Tspr18_2_V_1>>32'sd51))))  begin if ((xpc10==10'sd415/*415:xpc10*/)) 
                   begin 
                           xpc10 <= 10'sd416/*416:xpc10*/;
                           Tsf0SPILL12_256 <= rtl_sign_extend6((32'sd0/*0:USA146*/==(32'sd0/*0:USA144*/==(64'sh7_ffff_ffff_ffff&Tspr18_2_V_1
                          ))));

                           end 
                           end 
                   else if ((xpc10==10'sd415/*415:xpc10*/))  begin 
                           xpc10 <= 10'sd421/*421:xpc10*/;
                           Tspr18_2_V_4 <= 1'h0;
                           Tsf0SPILL12_256 <= 32'sd0;
                           end 
                          if ((32'sd4094/*4094:USA136*/==(64'shfff&(Tspr18_2_V_0>>32'sd51))))  begin if ((xpc10==10'sd413/*413:xpc10*/)) 
                   begin 
                           xpc10 <= 10'sd414/*414:xpc10*/;
                           Tsf0SPILL10_256 <= rtl_sign_extend6((32'sd0/*0:USA140*/==(32'sd0/*0:USA138*/==(64'sh7_ffff_ffff_ffff&Tspr18_2_V_0
                          ))));

                           end 
                           end 
                   else if ((xpc10==10'sd413/*413:xpc10*/))  begin 
                           xpc10 <= 10'sd422/*422:xpc10*/;
                           Tspr18_2_V_2 <= 1'h0;
                           Tsf0SPILL10_256 <= 32'sd0;
                           end 
                          if ((xpc10==10'sd358/*358:xpc10*/))  begin 
                      if (!Tspr27_2_V_2 && !Tspr27_2_V_4 && !Tspr27_2_V_3)  begin 
                               xpc10 <= 10'sd360/*360:xpc10*/;
                               Tss2_SPILL_256 <= Tspr27_2_V_0;
                               end 
                              if (!Tspr27_2_V_2 && !Tspr27_2_V_4 && Tspr27_2_V_3)  begin 
                               xpc10 <= 10'sd360/*360:xpc10*/;
                               Tss2_SPILL_256 <= Tspr27_2_V_1;
                               end 
                              if (Tspr27_2_V_2 || Tspr27_2_V_4)  begin if (Tspr27_2_V_2 || Tspr27_2_V_4)  xpc10 <= 10'sd359/*359:xpc10*/;
                               end 
                           end 
                      if ((32'sd4094/*4094:USA128*/==(64'shfff&(Tspr27_2_V_1>>32'sd51))))  begin if ((xpc10==10'sd355/*355:xpc10*/)) 
                   begin 
                           xpc10 <= 10'sd356/*356:xpc10*/;
                           Tsf0SPILL12_256 <= rtl_sign_extend6((32'sd0/*0:USA132*/==(32'sd0/*0:USA130*/==(64'sh7_ffff_ffff_ffff&Tspr27_2_V_1
                          ))));

                           end 
                           end 
                   else if ((xpc10==10'sd355/*355:xpc10*/))  begin 
                           xpc10 <= 10'sd361/*361:xpc10*/;
                           Tspr27_2_V_4 <= 1'h0;
                           Tsf0SPILL12_256 <= 32'sd0;
                           end 
                          if ((32'sd4094/*4094:USA122*/==(64'shfff&(Tspr27_2_V_0>>32'sd51))))  begin if ((xpc10==10'sd353/*353:xpc10*/)) 
                   begin 
                           xpc10 <= 10'sd354/*354:xpc10*/;
                           Tsf0SPILL10_256 <= rtl_sign_extend6((32'sd0/*0:USA126*/==(32'sd0/*0:USA124*/==(64'sh7_ffff_ffff_ffff&Tspr27_2_V_0
                          ))));

                           end 
                           end 
                   else if ((xpc10==10'sd353/*353:xpc10*/))  begin 
                           xpc10 <= 10'sd362/*362:xpc10*/;
                           Tspr27_2_V_2 <= 1'h0;
                           Tsf0SPILL10_256 <= 32'sd0;
                           end 
                          if ((xpc10==10'sd335/*335:xpc10*/))  begin 
                      if (!Tspr21_3_V_2 && !Tspr21_3_V_4 && !Tspr21_3_V_3)  begin 
                               xpc10 <= 10'sd337/*337:xpc10*/;
                               Tsa1_SPILL_256 <= Tspr21_3_V_0;
                               end 
                              if (!Tspr21_3_V_2 && !Tspr21_3_V_4 && Tspr21_3_V_3)  begin 
                               xpc10 <= 10'sd337/*337:xpc10*/;
                               Tsa1_SPILL_256 <= Tspr21_3_V_1;
                               end 
                              if (Tspr21_3_V_2 || Tspr21_3_V_4)  begin if (Tspr21_3_V_2 || Tspr21_3_V_4)  xpc10 <= 10'sd336/*336:xpc10*/;
                               end 
                           end 
                      if ((32'sd4094/*4094:USA112*/==(64'shfff&(Tspr21_3_V_1>>32'sd51))))  begin if ((xpc10==10'sd332/*332:xpc10*/)) 
                   begin 
                           xpc10 <= 10'sd333/*333:xpc10*/;
                           Tsf0SPILL12_256 <= rtl_sign_extend6((32'sd0/*0:USA116*/==(32'sd0/*0:USA114*/==(64'sh7_ffff_ffff_ffff&Tspr21_3_V_1
                          ))));

                           end 
                           end 
                   else if ((xpc10==10'sd332/*332:xpc10*/))  begin 
                           xpc10 <= 10'sd338/*338:xpc10*/;
                           Tspr21_3_V_4 <= 1'h0;
                           Tsf0SPILL12_256 <= 32'sd0;
                           end 
                          if ((32'sd4094/*4094:USA106*/==(64'shfff&(Tspr21_3_V_0>>32'sd51))))  begin if ((xpc10==10'sd330/*330:xpc10*/)) 
                   begin 
                           xpc10 <= 10'sd331/*331:xpc10*/;
                           Tsf0SPILL10_256 <= rtl_sign_extend6((32'sd0/*0:USA110*/==(32'sd0/*0:USA108*/==(64'sh7_ffff_ffff_ffff&Tspr21_3_V_0
                          ))));

                           end 
                           end 
                   else if ((xpc10==10'sd330/*330:xpc10*/))  begin 
                           xpc10 <= 10'sd339/*339:xpc10*/;
                           Tspr21_3_V_2 <= 1'h0;
                           Tsf0SPILL10_256 <= 32'sd0;
                           end 
                          if ((xpc10==10'sd314/*314:xpc10*/))  begin 
                      if (!Tspr12_2_V_2 && !Tspr12_2_V_4 && !Tspr12_2_V_3)  begin 
                               xpc10 <= 10'sd316/*316:xpc10*/;
                               Tsa1_SPILL_256 <= Tspr12_2_V_0;
                               end 
                              if (!Tspr12_2_V_2 && !Tspr12_2_V_4 && Tspr12_2_V_3)  begin 
                               xpc10 <= 10'sd316/*316:xpc10*/;
                               Tsa1_SPILL_256 <= Tspr12_2_V_1;
                               end 
                              if (Tspr12_2_V_2 || Tspr12_2_V_4)  begin if (Tspr12_2_V_2 || Tspr12_2_V_4)  xpc10 <= 10'sd315/*315:xpc10*/;
                               end 
                           end 
                      if ((32'sd4094/*4094:USA98*/==(64'shfff&(Tspr12_2_V_1>>32'sd51))))  begin if ((xpc10==10'sd311/*311:xpc10*/))  begin 
                           xpc10 <= 10'sd312/*312:xpc10*/;
                           Tsf0SPILL12_256 <= rtl_sign_extend6((32'sd0/*0:USA102*/==(32'sd0/*0:USA100*/==(64'sh7_ffff_ffff_ffff&Tspr12_2_V_1
                          ))));

                           end 
                           end 
                   else if ((xpc10==10'sd311/*311:xpc10*/))  begin 
                           xpc10 <= 10'sd317/*317:xpc10*/;
                           Tspr12_2_V_4 <= 1'h0;
                           Tsf0SPILL12_256 <= 32'sd0;
                           end 
                          if ((32'sd4094/*4094:USA92*/==(64'shfff&(Tspr12_2_V_0>>32'sd51))))  begin if ((xpc10==10'sd309/*309:xpc10*/)) 
                   begin 
                           xpc10 <= 10'sd310/*310:xpc10*/;
                           Tsf0SPILL10_256 <= rtl_sign_extend6((32'sd0/*0:USA96*/==(32'sd0/*0:USA94*/==(64'sh7_ffff_ffff_ffff&Tspr12_2_V_0
                          ))));

                           end 
                           end 
                   else if ((xpc10==10'sd309/*309:xpc10*/))  begin 
                           xpc10 <= 10'sd318/*318:xpc10*/;
                           Tspr12_2_V_2 <= 1'h0;
                           Tsf0SPILL10_256 <= 32'sd0;
                           end 
                          
              case (xpc10)
                  10'sd241/*241:xpc10*/:  begin 
                      if (!Tspr3_2_V_2 && !Tspr3_2_V_4 && !Tspr3_2_V_3)  begin 
                               xpc10 <= 10'sd243/*243:xpc10*/;
                               Tsa1_SPILL_256 <= Tspr3_2_V_0;
                               end 
                              if (!Tspr3_2_V_2 && !Tspr3_2_V_4 && Tspr3_2_V_3)  begin 
                               xpc10 <= 10'sd243/*243:xpc10*/;
                               Tsa1_SPILL_256 <= Tspr3_2_V_1;
                               end 
                              if (Tspr3_2_V_2 || Tspr3_2_V_4)  begin if (Tspr3_2_V_2 || Tspr3_2_V_4)  xpc10 <= 10'sd242/*242:xpc10*/;
                               end 
                           end 
                      
                  10'sd245/*245:xpc10*/:  begin 
                      if ((32'sd2047/*2047:USA166*/!=rtl_signed_bitextract9(64'sh7ff&((64'sh_7fff_ffff_ffff_ffff&Tdsi3_5_V_1)>>32'sd52
                      ))))  begin 
                               xpc10 <= 10'sd258/*258:xpc10*/;
                               Tsfl0_3_V_0 <= 1'h0;
                               end 
                              if ((32'sd2047/*2047:USA166*/==rtl_signed_bitextract9(64'sh7ff&((64'sh_7fff_ffff_ffff_ffff&Tdsi3_5_V_1)>>
                      32'sd52))) && (32'sd0/*0:USA168*/==(52'sd4503599627370495&Tdsi3_5_V_1)))  begin 
                               xpc10 <= 10'sd258/*258:xpc10*/;
                               Tsfl0_3_V_0 <= 1'h0;
                               end 
                              if ((32'sd2047/*2047:USA166*/==rtl_signed_bitextract9(64'sh7ff&((64'sh_7fff_ffff_ffff_ffff&Tdsi3_5_V_1)>>
                      32'sd52))) && (32'sd0/*0:USA168*/!=(52'sd4503599627370495&Tdsi3_5_V_1)))  xpc10 <= 10'sd246/*246:xpc10*/;
                           end 
                      
                  10'sd271/*271:xpc10*/: if (($signed(Tsad1_3_V_5)<64'sh0))  begin 
                           xpc10 <= 10'sd272/*272:xpc10*/;
                           Tsad1_3_V_5 <= Tsad1_3_V_3+Tsad1_3_V_4;
                           end 
                           else  begin 
                           xpc10 <= 10'sd274/*274:xpc10*/;
                           Tsro28_4_V_1 <= Tsad1_3_V_5;
                           Tsro28_4_V_0 <= rtl_signed_bitextract0(Tsad1_3_V_2);
                           end 
                          endcase
              if ((32'sd4094/*4094:USA84*/==(64'shfff&(Tspr3_2_V_1>>32'sd51))))  begin if ((xpc10==10'sd238/*238:xpc10*/))  begin 
                           xpc10 <= 10'sd239/*239:xpc10*/;
                           Tsf0SPILL12_256 <= rtl_sign_extend6((32'sd0/*0:USA88*/==(32'sd0/*0:USA86*/==(64'sh7_ffff_ffff_ffff&Tspr3_2_V_1
                          ))));

                           end 
                           end 
                   else if ((xpc10==10'sd238/*238:xpc10*/))  begin 
                           xpc10 <= 10'sd264/*264:xpc10*/;
                           Tspr3_2_V_4 <= 1'h0;
                           Tsf0SPILL12_256 <= 32'sd0;
                           end 
                          if ((32'sd4094/*4094:USA78*/==(64'shfff&(Tspr3_2_V_0>>32'sd51))))  begin if ((xpc10==10'sd236/*236:xpc10*/)) 
                   begin 
                           xpc10 <= 10'sd237/*237:xpc10*/;
                           Tsf0SPILL10_256 <= rtl_sign_extend6((32'sd0/*0:USA82*/==(32'sd0/*0:USA80*/==(64'sh7_ffff_ffff_ffff&Tspr3_2_V_0
                          ))));

                           end 
                           end 
                   else if ((xpc10==10'sd236/*236:xpc10*/))  begin 
                           xpc10 <= 10'sd265/*265:xpc10*/;
                           Tspr3_2_V_2 <= 1'h0;
                           Tsf0SPILL10_256 <= 32'sd0;
                           end 
                          if ((xpc10==10'sd224/*224:xpc10*/))  begin 
                      if (!Tspr2_2_V_2 && !Tspr2_2_V_4 && !Tspr2_2_V_3)  begin 
                               xpc10 <= 10'sd226/*226:xpc10*/;
                               Tsf1SPILL10_256 <= Tspr2_2_V_0;
                               end 
                              if (!Tspr2_2_V_2 && !Tspr2_2_V_4 && Tspr2_2_V_3)  begin 
                               xpc10 <= 10'sd226/*226:xpc10*/;
                               Tsf1SPILL10_256 <= Tspr2_2_V_1;
                               end 
                              if (Tspr2_2_V_2 || Tspr2_2_V_4)  begin if (Tspr2_2_V_2 || Tspr2_2_V_4)  xpc10 <= 10'sd225/*225:xpc10*/;
                               end 
                           end 
                      if ((32'sd4094/*4094:USA44*/==(64'shfff&(Tspr2_2_V_1>>32'sd51))))  begin if ((xpc10==10'sd221/*221:xpc10*/))  begin 
                           xpc10 <= 10'sd222/*222:xpc10*/;
                           Tsf0SPILL12_256 <= rtl_sign_extend6((32'sd0/*0:USA48*/==(32'sd0/*0:USA46*/==(64'sh7_ffff_ffff_ffff&Tspr2_2_V_1
                          ))));

                           end 
                           end 
                   else if ((xpc10==10'sd221/*221:xpc10*/))  begin 
                           xpc10 <= 10'sd451/*451:xpc10*/;
                           Tspr2_2_V_4 <= 1'h0;
                           Tsf0SPILL12_256 <= 32'sd0;
                           end 
                          if ((32'sd4094/*4094:USA38*/==(64'shfff&(Tspr2_2_V_0>>32'sd51))))  begin if ((xpc10==10'sd219/*219:xpc10*/)) 
                   begin 
                           xpc10 <= 10'sd220/*220:xpc10*/;
                           Tsf0SPILL10_256 <= rtl_sign_extend6((32'sd0/*0:USA42*/==(32'sd0/*0:USA40*/==(64'sh7_ffff_ffff_ffff&Tspr2_2_V_0
                          ))));

                           end 
                           end 
                   else if ((xpc10==10'sd219/*219:xpc10*/))  begin 
                           xpc10 <= 10'sd452/*452:xpc10*/;
                           Tspr2_2_V_2 <= 1'h0;
                           Tsf0SPILL10_256 <= 32'sd0;
                           end 
                          if ((Tspr4_3_V_2 || Tspr4_3_V_4) && (xpc10==10'sd209/*209:xpc10*/))  xpc10 <= 10'sd210/*210:xpc10*/;
                  if ((Tspr4_3_V_2 || Tspr4_3_V_4) && (xpc10==10'sd191/*191:xpc10*/))  xpc10 <= 10'sd192/*192:xpc10*/;
                  
              case (xpc10)
                  10'sd254/*254:xpc10*/:  begin 
                       xpc10 <= 10'sd255/*255:xpc10*/;
                       done <= 1'h1;
                       end 
                      
                  10'sd256/*256:xpc10*/:  begin 
                       xpc10 <= 10'sd255/*255:xpc10*/;
                       done <= 1'h1;
                       end 
                      
                  10'sd258/*258:xpc10*/: if ((64'sh0<((64'sh_7fff_ffff_ffff_ffff&Tdsi3_5_V_1)>>32'sd63)))  begin 
                           xpc10 <= 10'sd259/*259:xpc10*/;
                           Tsfl0_3_V_1 <= 1'h1;
                           end 
                           else  begin 
                           xpc10 <= 10'sd259/*259:xpc10*/;
                           Tsfl0_3_V_1 <= 1'h0;
                           end 
                          
                  10'sd277/*277:xpc10*/: if (Tsfl1_22_V_0)  begin 
                           xpc10 <= 10'sd278/*278:xpc10*/;
                           fastspilldup64 <= 64'h_fff0_0000_0000_0000;
                           end 
                           else  begin 
                           xpc10 <= 10'sd278/*278:xpc10*/;
                           fastspilldup64 <= 64'h_7ff0_0000_0000_0000;
                           end 
                          
                  10'sd381/*381:xpc10*/: if (Tssu2_4_V_0)  begin 
                           xpc10 <= 10'sd382/*382:xpc10*/;
                           fastspilldup72 <= 64'h_fff0_0000_0000_0000;
                           end 
                           else  begin 
                           xpc10 <= 10'sd382/*382:xpc10*/;
                           fastspilldup72 <= 64'h_7ff0_0000_0000_0000;
                           end 
                          
                  10'sd507/*507:xpc10*/: if ((Tsfl1_18_V_6<Tsfl1_18_V_7))  begin 
                           xpc10 <= 10'sd574/*574:xpc10*/;
                           Tses25_5_V_0 <= (Tsfl1_18_V_7>>32'sd32);
                           end 
                           else  begin 
                           xpc10 <= 10'sd508/*508:xpc10*/;
                           Tsfl1_18_V_8 <= 64'h_ffff_ffff_ffff_ffff;
                           end 
                          
                  10'sd622/*622:xpc10*/: if ((Tsco5_4_V_0<32'sh100_0000))  begin 
                           xpc10 <= 10'sd623/*623:xpc10*/;
                           Tsco5_4_V_1 <= rtl_unsigned_bitextract3(8'd8+Tsco5_4_V_1);
                           end 
                           else  begin 
                           xpc10 <= 10'sd625/*625:xpc10*/;
                           Tsco5_4_V_1 <= rtl_unsigned_bitextract3(Tsco5_4_V_1+A_8_US_CC_SCALbx14_ARA0[$unsigned((Tsco5_4_V_0>>32'sd24
                          ))]);

                           end 
                          
                  10'sd700/*700:xpc10*/: if (Tsfl1_7_V_2)  begin 
                           xpc10 <= 10'sd701/*701:xpc10*/;
                           fastspilldup32 <= 64'h_fff0_0000_0000_0000;
                           end 
                           else  begin 
                           xpc10 <= 10'sd701/*701:xpc10*/;
                           fastspilldup32 <= 64'h_7ff0_0000_0000_0000;
                           end 
                          
                  10'sd798/*798:xpc10*/: if (Tsfl0_9_V_2)  begin 
                           xpc10 <= 10'sd799/*799:xpc10*/;
                           fastspilldup22 <= 64'h_fff0_0000_0000_0000;
                           end 
                           else  begin 
                           xpc10 <= 10'sd799/*799:xpc10*/;
                           fastspilldup22 <= 64'h_7ff0_0000_0000_0000;
                           end 
                          endcase
              if ((32'sd0/*0:USA176*/==(Tdbm0_3_V_2^A_64_US_CC_SCALbx10_ARA0[Tdbm0_3_V_1])))  begin if ((xpc10==10'sd251/*251:xpc10*/)) 
                   begin 
                           xpc10 <= 10'sd253/*253:xpc10*/;
                           Tdbm0_3_V_1 <= 32'sd1+Tdbm0_3_V_1;
                           end 
                           end 
                   else if ((xpc10==10'sd251/*251:xpc10*/))  xpc10 <= 10'sd252/*252:xpc10*/;
                      
              case (xpc10)
                  10'sd0/*0:xpc10*/:  begin 
                       xpc10 <= 10'sd1/*1:xpc10*/;
                       dfsin_gloops <= 32'sd0;
                       end 
                      
                  10'sd1/*1:xpc10*/:  begin 
                       xpc10 <= 10'sd2/*2:xpc10*/;
                       A_64_US_CC_SCALbx12_ARB0[64'd0] <= 64'd0;
                       end 
                      
                  10'sd2/*2:xpc10*/:  begin 
                       xpc10 <= 10'sd3/*3:xpc10*/;
                       A_64_US_CC_SCALbx12_ARB0[64'd2] <= 64'sh_3fd6_5717_fced_55c1;
                       A_64_US_CC_SCALbx12_ARB0[64'd1] <= 64'sh_3fc6_5717_fced_55c1;
                       end 
                      
                  10'sd3/*3:xpc10*/:  begin 
                       xpc10 <= 10'sd4/*4:xpc10*/;
                       A_64_US_CC_SCALbx12_ARB0[64'd4] <= 64'sh_3fe6_5717_fced_55c1;
                       A_64_US_CC_SCALbx12_ARB0[64'd3] <= 64'sh_3fe0_c151_fdb2_0051;
                       end 
                      
                  10'sd4/*4:xpc10*/:  begin 
                       xpc10 <= 10'sd5/*5:xpc10*/;
                       A_64_US_CC_SCALbx12_ARB0[64'd6] <= 64'sh_3ff0_c151_fdb2_0051;
                       A_64_US_CC_SCALbx12_ARB0[64'd5] <= 64'sh_3feb_ecdd_fc28_ab31;
                       end 
                      
                  10'sd5/*5:xpc10*/:  begin 
                       xpc10 <= 10'sd6/*6:xpc10*/;
                       A_64_US_CC_SCALbx12_ARB0[64'd8] <= 64'sh_3ff6_5717_fced_55c1;
                       A_64_US_CC_SCALbx12_ARB0[64'd7] <= 64'sh_3ff3_8c34_fd4f_ab09;
                       end 
                      
                  10'sd6/*6:xpc10*/:  begin 
                       xpc10 <= 10'sd7/*7:xpc10*/;
                       A_64_US_CC_SCALbx12_ARB0[64'd10] <= 64'sh_3ffb_ecdd_fc28_ab31;
                       A_64_US_CC_SCALbx12_ARB0[64'd9] <= 64'sh_3ff9_21fa_fc8b_0079;
                       end 
                      
                  10'sd7/*7:xpc10*/:  begin 
                       xpc10 <= 10'sd8/*8:xpc10*/;
                       A_64_US_CC_SCALbx12_ARB0[64'd12] <= 64'sh_4000_c151_fdb2_0051;
                       A_64_US_CC_SCALbx12_ARB0[64'd11] <= 64'sh_3ffe_b7c0_fbc6_55e9;
                       end 
                      
                  10'sd8/*8:xpc10*/:  begin 
                       xpc10 <= 10'sd9/*9:xpc10*/;
                       A_64_US_CC_SCALbx12_ARB0[64'd14] <= 64'sh_4003_8c34_fd4f_ab09;
                       A_64_US_CC_SCALbx12_ARB0[64'd13] <= 64'sh_4002_26c3_7d80_d5ad;
                       end 
                      
                  10'sd9/*9:xpc10*/:  begin 
                       xpc10 <= 10'sd10/*10:xpc10*/;
                       A_64_US_CC_SCALbx12_ARB0[64'd16] <= 64'sh_4006_5717_fced_55c1;
                       A_64_US_CC_SCALbx12_ARB0[64'd15] <= 64'sh_4004_f1a6_7d1e_8065;
                       end 
                      
                  10'sd10/*10:xpc10*/:  begin 
                       xpc10 <= 10'sd11/*11:xpc10*/;
                       A_64_US_CC_SCALbx12_ARB0[64'd18] <= 64'sh_4009_21fa_fc8b_0079;
                       A_64_US_CC_SCALbx12_ARB0[64'd17] <= 64'sh_4007_bc89_7cbc_2b1d;
                       end 
                      
                  10'sd11/*11:xpc10*/:  begin 
                       xpc10 <= 10'sd12/*12:xpc10*/;
                       A_64_US_CC_SCALbx12_ARB0[64'd20] <= 64'sh_400b_ecdd_fc28_ab31;
                       A_64_US_CC_SCALbx12_ARB0[64'd19] <= 64'sh_400a_876c_7c59_d5d5;
                       end 
                      
                  10'sd12/*12:xpc10*/:  begin 
                       xpc10 <= 10'sd13/*13:xpc10*/;
                       A_64_US_CC_SCALbx12_ARB0[64'd22] <= 64'sh_400e_b7c0_fbc6_55e9;
                       A_64_US_CC_SCALbx12_ARB0[64'd21] <= 64'sh_400d_524f_7bf7_808d;
                       end 
                      
                  10'sd13/*13:xpc10*/:  begin 
                       xpc10 <= 10'sd14/*14:xpc10*/;
                       A_64_US_CC_SCALbx12_ARB0[64'd24] <= 64'sh_4010_c151_fdb2_0051;
                       A_64_US_CC_SCALbx12_ARB0[64'd23] <= 64'sh_4010_0e99_3dca_95a3;
                       end 
                      
                  10'sd14/*14:xpc10*/:  begin 
                       xpc10 <= 10'sd15/*15:xpc10*/;
                       A_64_US_CC_SCALbx12_ARB0[64'd26] <= 64'sh_4012_26c3_7d80_d5ad;
                       A_64_US_CC_SCALbx12_ARB0[64'd25] <= 64'sh_4011_740a_bd99_6aff;
                       end 
                      
                  10'sd15/*15:xpc10*/:  begin 
                       xpc10 <= 10'sd16/*16:xpc10*/;
                       A_64_US_CC_SCALbx12_ARB0[64'd28] <= 64'sh_4013_8c34_fd4f_ab09;
                       A_64_US_CC_SCALbx12_ARB0[64'd27] <= 64'sh_4012_d97c_3d68_405b;
                       end 
                      
                  10'sd16/*16:xpc10*/:  begin 
                       xpc10 <= 10'sd17/*17:xpc10*/;
                       A_64_US_CC_SCALbx12_ARB0[64'd30] <= 64'sh_4014_f1a6_7d1e_8065;
                       A_64_US_CC_SCALbx12_ARB0[64'd29] <= 64'sh_4014_3eed_bd37_15b7;
                       end 
                      
                  10'sd17/*17:xpc10*/:  begin 
                       xpc10 <= 10'sd18/*18:xpc10*/;
                       A_64_US_CC_SCALbx12_ARB0[64'd32] <= 64'sh_4016_5717_fced_55c1;
                       A_64_US_CC_SCALbx12_ARB0[64'd31] <= 64'sh_4015_a45f_3d05_eb13;
                       end 
                      
                  10'sd18/*18:xpc10*/:  begin 
                       xpc10 <= 10'sd19/*19:xpc10*/;
                       A_64_US_CC_SCALbx12_ARB0[64'd34] <= 64'sh_4017_bc89_7cbc_2b1d;
                       A_64_US_CC_SCALbx12_ARB0[64'd33] <= 64'sh_4017_09d0_bcd4_c06f;
                       end 
                      
                  10'sd19/*19:xpc10*/:  begin 
                       xpc10 <= 10'sd20/*20:xpc10*/;
                       A_64_US_CC_SCALbx12_ARB0[64'd35] <= 64'sh_4018_6f42_3ca3_95cb;
                       end 
                      
                  10'sd21/*21:xpc10*/:  begin 
                       xpc10 <= 10'sd22/*22:xpc10*/;
                       A_64_US_CC_SCALbx10_ARA0[64'd1] <= 64'sh_3fc6_3a1a_335a_adcd;
                       A_64_US_CC_SCALbx10_ARA0[64'd0] <= 64'd0;
                       end 
                      
                  10'sd22/*22:xpc10*/:  begin 
                       xpc10 <= 10'sd23/*23:xpc10*/;
                       A_64_US_CC_SCALbx10_ARA0[64'd3] <= 64'sh_3fdf_ffff_91f9_aa91;
                       A_64_US_CC_SCALbx10_ARA0[64'd2] <= 64'sh_3fd5_e3a8_2b09_bf3e;
                       end 
                      
                  10'sd23/*23:xpc10*/:  begin 
                       xpc10 <= 10'sd24/*24:xpc10*/;
                       A_64_US_CC_SCALbx10_ARA0[64'd5] <= 64'sh_3fe8_836f_6726_14a6;
                       A_64_US_CC_SCALbx10_ARA0[64'd4] <= 64'sh_3fe4_91b7_16c2_42e3;
                       end 
                      
                  10'sd24/*24:xpc10*/:  begin 
                       xpc10 <= 10'sd25/*25:xpc10*/;
                       A_64_US_CC_SCALbx10_ARA0[64'd7] <= 64'sh_3fee_11f6_127e_28ad;
                       A_64_US_CC_SCALbx10_ARA0[64'd6] <= 64'sh_3feb_b67a_c40b_2bed;
                       end 
                      
                  10'sd25/*25:xpc10*/:  begin 
                       xpc10 <= 10'sd26/*26:xpc10*/;
                       A_64_US_CC_SCALbx10_ARA0[64'd9] <= 64'sh_3fef_ffff_e1cb_d7aa;
                       A_64_US_CC_SCALbx10_ARA0[64'd8] <= 64'sh_3fef_838b_6adf_fac0;
                       end 
                      
                  10'sd26/*26:xpc10*/:  begin 
                       xpc10 <= 10'sd27/*27:xpc10*/;
                       A_64_US_CC_SCALbx10_ARA0[64'd11] <= 64'sh_3fee_11f6_92d9_62b4;
                       A_64_US_CC_SCALbx10_ARA0[64'd10] <= 64'sh_3fef_838b_b014_7989;
                       end 
                      
                  10'sd27/*27:xpc10*/:  begin 
                       xpc10 <= 10'sd28/*28:xpc10*/;
                       A_64_US_CC_SCALbx10_ARA0[64'd13] <= 64'sh_3fe8_8370_9d4e_a869;
                       A_64_US_CC_SCALbx10_ARA0[64'd12] <= 64'sh_3feb_b67b_77c0_142d;
                       end 
                      
                  10'sd28/*28:xpc10*/:  begin 
                       xpc10 <= 10'sd29/*29:xpc10*/;
                       A_64_US_CC_SCALbx10_ARA0[64'd15] <= 64'sh_3fe0_0000_ea5f_43c8;
                       A_64_US_CC_SCALbx10_ARA0[64'd14] <= 64'sh_3fe4_91b8_1d72_d8e8;
                       end 
                      
                  10'sd29/*29:xpc10*/:  begin 
                       xpc10 <= 10'sd30/*30:xpc10*/;
                       A_64_US_CC_SCALbx10_ARA0[64'd17] <= 64'sh_3fc6_3a1d_2189_552c;
                       A_64_US_CC_SCALbx10_ARA0[64'd16] <= 64'sh_3fd5_e3aa_4e05_90c5;
                       end 
                      
                  10'sd30/*30:xpc10*/:  begin 
                       xpc10 <= 10'sd31/*31:xpc10*/;
                       A_64_US_CC_SCALbx10_ARA0[64'd19] <= -64'sh_4039_c5eb_bb22_4c84;
                       A_64_US_CC_SCALbx10_ARA0[64'd18] <= 64'sh_3ea6_aedf_fc45_4b91;
                       end 
                      
                  10'sd31/*31:xpc10*/:  begin 
                       xpc10 <= 10'sd32/*32:xpc10*/;
                       A_64_US_CC_SCALbx10_ARA0[64'd21] <= -64'sh_4020_0002_b6b3_0695;
                       A_64_US_CC_SCALbx10_ARA0[64'd20] <= -64'sh_402a_1c5b_1970_70c2;
                       end 
                      
                  10'sd32/*32:xpc10*/:  begin 
                       xpc10 <= 10'sd33/*33:xpc10*/;
                       A_64_US_CC_SCALbx10_ARA0[64'd23] <= -64'sh_4017_7c91_4d23_07eb;
                       A_64_US_CC_SCALbx10_ARA0[64'd22] <= -64'sh_401b_6e49_e346_5c2d;
                       end 
                      
                  10'sd33/*33:xpc10*/:  begin 
                       xpc10 <= 10'sd34/*34:xpc10*/;
                       A_64_US_CC_SCALbx10_ARA0[64'd25] <= -64'sh_4011_ee0a_6ed2_dea9;
                       A_64_US_CC_SCALbx10_ARA0[64'd24] <= -64'sh_4014_4985_8bf5_51ce;
                       end 
                      
                  10'sd34/*34:xpc10*/:  begin 
                       xpc10 <= 10'sd35/*35:xpc10*/;
                       A_64_US_CC_SCALbx10_ARA0[64'd27] <= -64'sh_4010_0000_3d1a_2371;
                       A_64_US_CC_SCALbx10_ARA0[64'd26] <= -64'sh_4010_7c74_e539_b504;
                       end 
                      
                  10'sd35/*35:xpc10*/:  begin 
                       xpc10 <= 10'sd36/*36:xpc10*/;
                       A_64_US_CC_SCALbx10_ARA0[64'd29] <= -64'sh_4011_ee08_eed2_51d9;
                       A_64_US_CC_SCALbx10_ARA0[64'd28] <= -64'sh_4010_7c74_a15d_1816;
                       end 
                      
                  10'sd36/*36:xpc10*/:  begin 
                       xpc10 <= 10'sd37/*37:xpc10*/;
                       A_64_US_CC_SCALbx10_ARA0[64'd31] <= -64'sh_4017_7c8e_9190_287f;
                       A_64_US_CC_SCALbx10_ARA0[64'd30] <= -64'sh_4014_4983_d3ce_34b6;
                       end 
                      
                  10'sd37/*37:xpc10*/:  begin 
                       xpc10 <= 10'sd38/*38:xpc10*/;
                       A_64_US_CC_SCALbx10_ARA0[64'd33] <= -64'sh_401f_fffd_e2f3_5cf3;
                       A_64_US_CC_SCALbx10_ARA0[64'd32] <= -64'sh_401b_6e46_32e4_a2aa;
                       end 
                      
                  10'sd38/*38:xpc10*/:  begin 
                       xpc10 <= 10'sd39/*39:xpc10*/;
                       A_64_US_CC_SCALbx10_ARA0[64'd35] <= -64'sh_4039_c5dc_3b77_9c23;
                       A_64_US_CC_SCALbx10_ARA0[64'd34] <= -64'sh_402a_1c52_f596_3509;
                       end 
                      
                  10'sd39/*39:xpc10*/:  begin 
                       xpc10 <= 10'sd40/*40:xpc10*/;
                       done <= 1'h0;
                       end 
                      
                  10'sd41/*41:xpc10*/:  begin 
                       xpc10 <= 10'sd42/*42:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[32'd0] <= 8'h8;
                       end 
                      
                  10'sd42/*42:xpc10*/:  begin 
                       xpc10 <= 10'sd43/*43:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh2] <= 8'h6;
                       A_8_US_CC_SCALbx14_ARA0[64'sh1] <= 8'h7;
                       end 
                      
                  10'sd43/*43:xpc10*/:  begin 
                       xpc10 <= 10'sd44/*44:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh4] <= 8'h5;
                       A_8_US_CC_SCALbx14_ARA0[64'sh3] <= 8'h6;
                       end 
                      
                  10'sd44/*44:xpc10*/:  begin 
                       xpc10 <= 10'sd45/*45:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh6] <= 8'h5;
                       A_8_US_CC_SCALbx14_ARA0[64'sh5] <= 8'h5;
                       end 
                      
                  10'sd45/*45:xpc10*/:  begin 
                       xpc10 <= 10'sd46/*46:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh8] <= 8'h4;
                       A_8_US_CC_SCALbx14_ARA0[64'sh7] <= 8'h5;
                       end 
                      
                  10'sd46/*46:xpc10*/:  begin 
                       xpc10 <= 10'sd47/*47:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sha] <= 8'h4;
                       A_8_US_CC_SCALbx14_ARA0[64'sh9] <= 8'h4;
                       end 
                      
                  10'sd47/*47:xpc10*/:  begin 
                       xpc10 <= 10'sd48/*48:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'shc] <= 8'h4;
                       A_8_US_CC_SCALbx14_ARA0[64'shb] <= 8'h4;
                       end 
                      
                  10'sd48/*48:xpc10*/:  begin 
                       xpc10 <= 10'sd49/*49:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'she] <= 8'h4;
                       A_8_US_CC_SCALbx14_ARA0[64'shd] <= 8'h4;
                       end 
                      
                  10'sd49/*49:xpc10*/:  begin 
                       xpc10 <= 10'sd50/*50:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh10] <= 8'h3;
                       A_8_US_CC_SCALbx14_ARA0[64'shf] <= 8'h4;
                       end 
                      
                  10'sd50/*50:xpc10*/:  begin 
                       xpc10 <= 10'sd51/*51:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh12] <= 8'h3;
                       A_8_US_CC_SCALbx14_ARA0[64'sh11] <= 8'h3;
                       end 
                      
                  10'sd51/*51:xpc10*/:  begin 
                       xpc10 <= 10'sd52/*52:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh14] <= 8'h3;
                       A_8_US_CC_SCALbx14_ARA0[64'sh13] <= 8'h3;
                       end 
                      
                  10'sd52/*52:xpc10*/:  begin 
                       xpc10 <= 10'sd53/*53:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh16] <= 8'h3;
                       A_8_US_CC_SCALbx14_ARA0[64'sh15] <= 8'h3;
                       end 
                      
                  10'sd53/*53:xpc10*/:  begin 
                       xpc10 <= 10'sd54/*54:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh18] <= 8'h3;
                       A_8_US_CC_SCALbx14_ARA0[64'sh17] <= 8'h3;
                       end 
                      
                  10'sd54/*54:xpc10*/:  begin 
                       xpc10 <= 10'sd55/*55:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh1a] <= 8'h3;
                       A_8_US_CC_SCALbx14_ARA0[64'sh19] <= 8'h3;
                       end 
                      
                  10'sd55/*55:xpc10*/:  begin 
                       xpc10 <= 10'sd56/*56:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh1c] <= 8'h3;
                       A_8_US_CC_SCALbx14_ARA0[64'sh1b] <= 8'h3;
                       end 
                      
                  10'sd56/*56:xpc10*/:  begin 
                       xpc10 <= 10'sd57/*57:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh1e] <= 8'h3;
                       A_8_US_CC_SCALbx14_ARA0[64'sh1d] <= 8'h3;
                       end 
                      
                  10'sd57/*57:xpc10*/:  begin 
                       xpc10 <= 10'sd58/*58:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh20] <= 8'h2;
                       A_8_US_CC_SCALbx14_ARA0[64'sh1f] <= 8'h3;
                       end 
                      
                  10'sd58/*58:xpc10*/:  begin 
                       xpc10 <= 10'sd59/*59:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh22] <= 8'h2;
                       A_8_US_CC_SCALbx14_ARA0[64'sh21] <= 8'h2;
                       end 
                      
                  10'sd59/*59:xpc10*/:  begin 
                       xpc10 <= 10'sd60/*60:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh24] <= 8'h2;
                       A_8_US_CC_SCALbx14_ARA0[64'sh23] <= 8'h2;
                       end 
                      
                  10'sd60/*60:xpc10*/:  begin 
                       xpc10 <= 10'sd61/*61:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh26] <= 8'h2;
                       A_8_US_CC_SCALbx14_ARA0[64'sh25] <= 8'h2;
                       end 
                      
                  10'sd61/*61:xpc10*/:  begin 
                       xpc10 <= 10'sd62/*62:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh28] <= 8'h2;
                       A_8_US_CC_SCALbx14_ARA0[64'sh27] <= 8'h2;
                       end 
                      
                  10'sd62/*62:xpc10*/:  begin 
                       xpc10 <= 10'sd63/*63:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh2a] <= 8'h2;
                       A_8_US_CC_SCALbx14_ARA0[64'sh29] <= 8'h2;
                       end 
                      
                  10'sd63/*63:xpc10*/:  begin 
                       xpc10 <= 10'sd64/*64:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh2c] <= 8'h2;
                       A_8_US_CC_SCALbx14_ARA0[64'sh2b] <= 8'h2;
                       end 
                      
                  10'sd64/*64:xpc10*/:  begin 
                       xpc10 <= 10'sd65/*65:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh2e] <= 8'h2;
                       A_8_US_CC_SCALbx14_ARA0[64'sh2d] <= 8'h2;
                       end 
                      
                  10'sd65/*65:xpc10*/:  begin 
                       xpc10 <= 10'sd66/*66:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh30] <= 8'h2;
                       A_8_US_CC_SCALbx14_ARA0[64'sh2f] <= 8'h2;
                       end 
                      
                  10'sd66/*66:xpc10*/:  begin 
                       xpc10 <= 10'sd67/*67:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh32] <= 8'h2;
                       A_8_US_CC_SCALbx14_ARA0[64'sh31] <= 8'h2;
                       end 
                      
                  10'sd67/*67:xpc10*/:  begin 
                       xpc10 <= 10'sd68/*68:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh34] <= 8'h2;
                       A_8_US_CC_SCALbx14_ARA0[64'sh33] <= 8'h2;
                       end 
                      
                  10'sd68/*68:xpc10*/:  begin 
                       xpc10 <= 10'sd69/*69:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh36] <= 8'h2;
                       A_8_US_CC_SCALbx14_ARA0[64'sh35] <= 8'h2;
                       end 
                      
                  10'sd69/*69:xpc10*/:  begin 
                       xpc10 <= 10'sd70/*70:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh38] <= 8'h2;
                       A_8_US_CC_SCALbx14_ARA0[64'sh37] <= 8'h2;
                       end 
                      
                  10'sd70/*70:xpc10*/:  begin 
                       xpc10 <= 10'sd71/*71:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh3a] <= 8'h2;
                       A_8_US_CC_SCALbx14_ARA0[64'sh39] <= 8'h2;
                       end 
                      
                  10'sd71/*71:xpc10*/:  begin 
                       xpc10 <= 10'sd72/*72:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh3c] <= 8'h2;
                       A_8_US_CC_SCALbx14_ARA0[64'sh3b] <= 8'h2;
                       end 
                      
                  10'sd72/*72:xpc10*/:  begin 
                       xpc10 <= 10'sd73/*73:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh3e] <= 8'h2;
                       A_8_US_CC_SCALbx14_ARA0[64'sh3d] <= 8'h2;
                       end 
                      
                  10'sd73/*73:xpc10*/:  begin 
                       xpc10 <= 10'sd74/*74:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh40] <= 8'h1;
                       A_8_US_CC_SCALbx14_ARA0[64'sh3f] <= 8'h2;
                       end 
                      
                  10'sd74/*74:xpc10*/:  begin 
                       xpc10 <= 10'sd75/*75:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh42] <= 8'h1;
                       A_8_US_CC_SCALbx14_ARA0[64'sh41] <= 8'h1;
                       end 
                      
                  10'sd75/*75:xpc10*/:  begin 
                       xpc10 <= 10'sd76/*76:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh44] <= 8'h1;
                       A_8_US_CC_SCALbx14_ARA0[64'sh43] <= 8'h1;
                       end 
                      
                  10'sd76/*76:xpc10*/:  begin 
                       xpc10 <= 10'sd77/*77:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh46] <= 8'h1;
                       A_8_US_CC_SCALbx14_ARA0[64'sh45] <= 8'h1;
                       end 
                      
                  10'sd77/*77:xpc10*/:  begin 
                       xpc10 <= 10'sd78/*78:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh48] <= 8'h1;
                       A_8_US_CC_SCALbx14_ARA0[64'sh47] <= 8'h1;
                       end 
                      
                  10'sd78/*78:xpc10*/:  begin 
                       xpc10 <= 10'sd79/*79:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh4a] <= 8'h1;
                       A_8_US_CC_SCALbx14_ARA0[64'sh49] <= 8'h1;
                       end 
                      
                  10'sd79/*79:xpc10*/:  begin 
                       xpc10 <= 10'sd80/*80:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh4c] <= 8'h1;
                       A_8_US_CC_SCALbx14_ARA0[64'sh4b] <= 8'h1;
                       end 
                      
                  10'sd80/*80:xpc10*/:  begin 
                       xpc10 <= 10'sd81/*81:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh4e] <= 8'h1;
                       A_8_US_CC_SCALbx14_ARA0[64'sh4d] <= 8'h1;
                       end 
                      
                  10'sd81/*81:xpc10*/:  begin 
                       xpc10 <= 10'sd82/*82:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh50] <= 8'h1;
                       A_8_US_CC_SCALbx14_ARA0[64'sh4f] <= 8'h1;
                       end 
                      
                  10'sd82/*82:xpc10*/:  begin 
                       xpc10 <= 10'sd83/*83:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh52] <= 8'h1;
                       A_8_US_CC_SCALbx14_ARA0[64'sh51] <= 8'h1;
                       end 
                      
                  10'sd83/*83:xpc10*/:  begin 
                       xpc10 <= 10'sd84/*84:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh54] <= 8'h1;
                       A_8_US_CC_SCALbx14_ARA0[64'sh53] <= 8'h1;
                       end 
                      
                  10'sd84/*84:xpc10*/:  begin 
                       xpc10 <= 10'sd85/*85:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh56] <= 8'h1;
                       A_8_US_CC_SCALbx14_ARA0[64'sh55] <= 8'h1;
                       end 
                      
                  10'sd85/*85:xpc10*/:  begin 
                       xpc10 <= 10'sd86/*86:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh58] <= 8'h1;
                       A_8_US_CC_SCALbx14_ARA0[64'sh57] <= 8'h1;
                       end 
                      
                  10'sd86/*86:xpc10*/:  begin 
                       xpc10 <= 10'sd87/*87:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh5a] <= 8'h1;
                       A_8_US_CC_SCALbx14_ARA0[64'sh59] <= 8'h1;
                       end 
                      
                  10'sd87/*87:xpc10*/:  begin 
                       xpc10 <= 10'sd88/*88:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh5c] <= 8'h1;
                       A_8_US_CC_SCALbx14_ARA0[64'sh5b] <= 8'h1;
                       end 
                      
                  10'sd88/*88:xpc10*/:  begin 
                       xpc10 <= 10'sd89/*89:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh5e] <= 8'h1;
                       A_8_US_CC_SCALbx14_ARA0[64'sh5d] <= 8'h1;
                       end 
                      
                  10'sd89/*89:xpc10*/:  begin 
                       xpc10 <= 10'sd90/*90:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh60] <= 8'h1;
                       A_8_US_CC_SCALbx14_ARA0[64'sh5f] <= 8'h1;
                       end 
                      
                  10'sd90/*90:xpc10*/:  begin 
                       xpc10 <= 10'sd91/*91:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh62] <= 8'h1;
                       A_8_US_CC_SCALbx14_ARA0[64'sh61] <= 8'h1;
                       end 
                      
                  10'sd91/*91:xpc10*/:  begin 
                       xpc10 <= 10'sd92/*92:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh64] <= 8'h1;
                       A_8_US_CC_SCALbx14_ARA0[64'sh63] <= 8'h1;
                       end 
                      
                  10'sd92/*92:xpc10*/:  begin 
                       xpc10 <= 10'sd93/*93:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh66] <= 8'h1;
                       A_8_US_CC_SCALbx14_ARA0[64'sh65] <= 8'h1;
                       end 
                      
                  10'sd93/*93:xpc10*/:  begin 
                       xpc10 <= 10'sd94/*94:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh68] <= 8'h1;
                       A_8_US_CC_SCALbx14_ARA0[64'sh67] <= 8'h1;
                       end 
                      
                  10'sd94/*94:xpc10*/:  begin 
                       xpc10 <= 10'sd95/*95:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh6a] <= 8'h1;
                       A_8_US_CC_SCALbx14_ARA0[64'sh69] <= 8'h1;
                       end 
                      
                  10'sd95/*95:xpc10*/:  begin 
                       xpc10 <= 10'sd96/*96:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh6c] <= 8'h1;
                       A_8_US_CC_SCALbx14_ARA0[64'sh6b] <= 8'h1;
                       end 
                      
                  10'sd96/*96:xpc10*/:  begin 
                       xpc10 <= 10'sd97/*97:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh6e] <= 8'h1;
                       A_8_US_CC_SCALbx14_ARA0[64'sh6d] <= 8'h1;
                       end 
                      
                  10'sd97/*97:xpc10*/:  begin 
                       xpc10 <= 10'sd98/*98:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh70] <= 8'h1;
                       A_8_US_CC_SCALbx14_ARA0[64'sh6f] <= 8'h1;
                       end 
                      
                  10'sd98/*98:xpc10*/:  begin 
                       xpc10 <= 10'sd99/*99:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh72] <= 8'h1;
                       A_8_US_CC_SCALbx14_ARA0[64'sh71] <= 8'h1;
                       end 
                      
                  10'sd99/*99:xpc10*/:  begin 
                       xpc10 <= 10'sd100/*100:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh74] <= 8'h1;
                       A_8_US_CC_SCALbx14_ARA0[64'sh73] <= 8'h1;
                       end 
                      
                  10'sd100/*100:xpc10*/:  begin 
                       xpc10 <= 10'sd101/*101:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh76] <= 8'h1;
                       A_8_US_CC_SCALbx14_ARA0[64'sh75] <= 8'h1;
                       end 
                      
                  10'sd101/*101:xpc10*/:  begin 
                       xpc10 <= 10'sd102/*102:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh78] <= 8'h1;
                       A_8_US_CC_SCALbx14_ARA0[64'sh77] <= 8'h1;
                       end 
                      
                  10'sd102/*102:xpc10*/:  begin 
                       xpc10 <= 10'sd103/*103:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh7a] <= 8'h1;
                       A_8_US_CC_SCALbx14_ARA0[64'sh79] <= 8'h1;
                       end 
                      
                  10'sd103/*103:xpc10*/:  begin 
                       xpc10 <= 10'sd104/*104:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh7c] <= 8'h1;
                       A_8_US_CC_SCALbx14_ARA0[64'sh7b] <= 8'h1;
                       end 
                      
                  10'sd104/*104:xpc10*/:  begin 
                       xpc10 <= 10'sd105/*105:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh7e] <= 8'h1;
                       A_8_US_CC_SCALbx14_ARA0[64'sh7d] <= 8'h1;
                       end 
                      
                  10'sd105/*105:xpc10*/:  begin 
                       xpc10 <= 10'sd106/*106:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh80] <= 8'h0;
                       A_8_US_CC_SCALbx14_ARA0[64'sh7f] <= 8'h1;
                       end 
                      
                  10'sd106/*106:xpc10*/:  begin 
                       xpc10 <= 10'sd107/*107:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh82] <= 8'h0;
                       A_8_US_CC_SCALbx14_ARA0[64'sh81] <= 8'h0;
                       end 
                      
                  10'sd107/*107:xpc10*/:  begin 
                       xpc10 <= 10'sd108/*108:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh84] <= 8'h0;
                       A_8_US_CC_SCALbx14_ARA0[64'sh83] <= 8'h0;
                       end 
                      
                  10'sd108/*108:xpc10*/:  begin 
                       xpc10 <= 10'sd109/*109:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh86] <= 8'h0;
                       A_8_US_CC_SCALbx14_ARA0[64'sh85] <= 8'h0;
                       end 
                      
                  10'sd109/*109:xpc10*/:  begin 
                       xpc10 <= 10'sd110/*110:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh88] <= 8'h0;
                       A_8_US_CC_SCALbx14_ARA0[64'sh87] <= 8'h0;
                       end 
                      
                  10'sd110/*110:xpc10*/:  begin 
                       xpc10 <= 10'sd111/*111:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh8a] <= 8'h0;
                       A_8_US_CC_SCALbx14_ARA0[64'sh89] <= 8'h0;
                       end 
                      
                  10'sd111/*111:xpc10*/:  begin 
                       xpc10 <= 10'sd112/*112:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh8c] <= 8'h0;
                       A_8_US_CC_SCALbx14_ARA0[64'sh8b] <= 8'h0;
                       end 
                      
                  10'sd112/*112:xpc10*/:  begin 
                       xpc10 <= 10'sd113/*113:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh8e] <= 8'h0;
                       A_8_US_CC_SCALbx14_ARA0[64'sh8d] <= 8'h0;
                       end 
                      
                  10'sd113/*113:xpc10*/:  begin 
                       xpc10 <= 10'sd114/*114:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh90] <= 8'h0;
                       A_8_US_CC_SCALbx14_ARA0[64'sh8f] <= 8'h0;
                       end 
                      
                  10'sd114/*114:xpc10*/:  begin 
                       xpc10 <= 10'sd115/*115:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh92] <= 8'h0;
                       A_8_US_CC_SCALbx14_ARA0[64'sh91] <= 8'h0;
                       end 
                      
                  10'sd115/*115:xpc10*/:  begin 
                       xpc10 <= 10'sd116/*116:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh94] <= 8'h0;
                       A_8_US_CC_SCALbx14_ARA0[64'sh93] <= 8'h0;
                       end 
                      
                  10'sd116/*116:xpc10*/:  begin 
                       xpc10 <= 10'sd117/*117:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh96] <= 8'h0;
                       A_8_US_CC_SCALbx14_ARA0[64'sh95] <= 8'h0;
                       end 
                      
                  10'sd117/*117:xpc10*/:  begin 
                       xpc10 <= 10'sd118/*118:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh98] <= 8'h0;
                       A_8_US_CC_SCALbx14_ARA0[64'sh97] <= 8'h0;
                       end 
                      
                  10'sd118/*118:xpc10*/:  begin 
                       xpc10 <= 10'sd119/*119:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh9a] <= 8'h0;
                       A_8_US_CC_SCALbx14_ARA0[64'sh99] <= 8'h0;
                       end 
                      
                  10'sd119/*119:xpc10*/:  begin 
                       xpc10 <= 10'sd120/*120:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh9c] <= 8'h0;
                       A_8_US_CC_SCALbx14_ARA0[64'sh9b] <= 8'h0;
                       end 
                      
                  10'sd120/*120:xpc10*/:  begin 
                       xpc10 <= 10'sd121/*121:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sh9e] <= 8'h0;
                       A_8_US_CC_SCALbx14_ARA0[64'sh9d] <= 8'h0;
                       end 
                      
                  10'sd121/*121:xpc10*/:  begin 
                       xpc10 <= 10'sd122/*122:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sha0] <= 8'h0;
                       A_8_US_CC_SCALbx14_ARA0[64'sh9f] <= 8'h0;
                       end 
                      
                  10'sd122/*122:xpc10*/:  begin 
                       xpc10 <= 10'sd123/*123:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sha2] <= 8'h0;
                       A_8_US_CC_SCALbx14_ARA0[64'sha1] <= 8'h0;
                       end 
                      
                  10'sd123/*123:xpc10*/:  begin 
                       xpc10 <= 10'sd124/*124:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sha4] <= 8'h0;
                       A_8_US_CC_SCALbx14_ARA0[64'sha3] <= 8'h0;
                       end 
                      
                  10'sd124/*124:xpc10*/:  begin 
                       xpc10 <= 10'sd125/*125:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sha6] <= 8'h0;
                       A_8_US_CC_SCALbx14_ARA0[64'sha5] <= 8'h0;
                       end 
                      
                  10'sd125/*125:xpc10*/:  begin 
                       xpc10 <= 10'sd126/*126:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'sha8] <= 8'h0;
                       A_8_US_CC_SCALbx14_ARA0[64'sha7] <= 8'h0;
                       end 
                      
                  10'sd126/*126:xpc10*/:  begin 
                       xpc10 <= 10'sd127/*127:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'shaa] <= 8'h0;
                       A_8_US_CC_SCALbx14_ARA0[64'sha9] <= 8'h0;
                       end 
                      
                  10'sd127/*127:xpc10*/:  begin 
                       xpc10 <= 10'sd128/*128:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'shac] <= 8'h0;
                       A_8_US_CC_SCALbx14_ARA0[64'shab] <= 8'h0;
                       end 
                      
                  10'sd128/*128:xpc10*/:  begin 
                       xpc10 <= 10'sd129/*129:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'shae] <= 8'h0;
                       A_8_US_CC_SCALbx14_ARA0[64'shad] <= 8'h0;
                       end 
                      
                  10'sd129/*129:xpc10*/:  begin 
                       xpc10 <= 10'sd130/*130:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'shb0] <= 8'h0;
                       A_8_US_CC_SCALbx14_ARA0[64'shaf] <= 8'h0;
                       end 
                      
                  10'sd130/*130:xpc10*/:  begin 
                       xpc10 <= 10'sd131/*131:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'shb2] <= 8'h0;
                       A_8_US_CC_SCALbx14_ARA0[64'shb1] <= 8'h0;
                       end 
                      
                  10'sd131/*131:xpc10*/:  begin 
                       xpc10 <= 10'sd132/*132:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'shb4] <= 8'h0;
                       A_8_US_CC_SCALbx14_ARA0[64'shb3] <= 8'h0;
                       end 
                      
                  10'sd132/*132:xpc10*/:  begin 
                       xpc10 <= 10'sd133/*133:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'shb6] <= 8'h0;
                       A_8_US_CC_SCALbx14_ARA0[64'shb5] <= 8'h0;
                       end 
                      
                  10'sd133/*133:xpc10*/:  begin 
                       xpc10 <= 10'sd134/*134:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'shb8] <= 8'h0;
                       A_8_US_CC_SCALbx14_ARA0[64'shb7] <= 8'h0;
                       end 
                      
                  10'sd134/*134:xpc10*/:  begin 
                       xpc10 <= 10'sd135/*135:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'shba] <= 8'h0;
                       A_8_US_CC_SCALbx14_ARA0[64'shb9] <= 8'h0;
                       end 
                      
                  10'sd135/*135:xpc10*/:  begin 
                       xpc10 <= 10'sd136/*136:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'shbc] <= 8'h0;
                       A_8_US_CC_SCALbx14_ARA0[64'shbb] <= 8'h0;
                       end 
                      
                  10'sd136/*136:xpc10*/:  begin 
                       xpc10 <= 10'sd137/*137:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'shbe] <= 8'h0;
                       A_8_US_CC_SCALbx14_ARA0[64'shbd] <= 8'h0;
                       end 
                      
                  10'sd137/*137:xpc10*/:  begin 
                       xpc10 <= 10'sd138/*138:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'shc0] <= 8'h0;
                       A_8_US_CC_SCALbx14_ARA0[64'shbf] <= 8'h0;
                       end 
                      
                  10'sd138/*138:xpc10*/:  begin 
                       xpc10 <= 10'sd139/*139:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'shc2] <= 8'h0;
                       A_8_US_CC_SCALbx14_ARA0[64'shc1] <= 8'h0;
                       end 
                      
                  10'sd139/*139:xpc10*/:  begin 
                       xpc10 <= 10'sd140/*140:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'shc4] <= 8'h0;
                       A_8_US_CC_SCALbx14_ARA0[64'shc3] <= 8'h0;
                       end 
                      
                  10'sd140/*140:xpc10*/:  begin 
                       xpc10 <= 10'sd141/*141:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'shc6] <= 8'h0;
                       A_8_US_CC_SCALbx14_ARA0[64'shc5] <= 8'h0;
                       end 
                      
                  10'sd141/*141:xpc10*/:  begin 
                       xpc10 <= 10'sd142/*142:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'shc8] <= 8'h0;
                       A_8_US_CC_SCALbx14_ARA0[64'shc7] <= 8'h0;
                       end 
                      
                  10'sd142/*142:xpc10*/:  begin 
                       xpc10 <= 10'sd143/*143:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'shca] <= 8'h0;
                       A_8_US_CC_SCALbx14_ARA0[64'shc9] <= 8'h0;
                       end 
                      
                  10'sd143/*143:xpc10*/:  begin 
                       xpc10 <= 10'sd144/*144:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'shcc] <= 8'h0;
                       A_8_US_CC_SCALbx14_ARA0[64'shcb] <= 8'h0;
                       end 
                      
                  10'sd144/*144:xpc10*/:  begin 
                       xpc10 <= 10'sd145/*145:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'shce] <= 8'h0;
                       A_8_US_CC_SCALbx14_ARA0[64'shcd] <= 8'h0;
                       end 
                      
                  10'sd145/*145:xpc10*/:  begin 
                       xpc10 <= 10'sd146/*146:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'shd0] <= 8'h0;
                       A_8_US_CC_SCALbx14_ARA0[64'shcf] <= 8'h0;
                       end 
                      
                  10'sd146/*146:xpc10*/:  begin 
                       xpc10 <= 10'sd147/*147:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'shd2] <= 8'h0;
                       A_8_US_CC_SCALbx14_ARA0[64'shd1] <= 8'h0;
                       end 
                      
                  10'sd147/*147:xpc10*/:  begin 
                       xpc10 <= 10'sd148/*148:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'shd4] <= 8'h0;
                       A_8_US_CC_SCALbx14_ARA0[64'shd3] <= 8'h0;
                       end 
                      
                  10'sd148/*148:xpc10*/:  begin 
                       xpc10 <= 10'sd149/*149:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'shd6] <= 8'h0;
                       A_8_US_CC_SCALbx14_ARA0[64'shd5] <= 8'h0;
                       end 
                      
                  10'sd149/*149:xpc10*/:  begin 
                       xpc10 <= 10'sd150/*150:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'shd8] <= 8'h0;
                       A_8_US_CC_SCALbx14_ARA0[64'shd7] <= 8'h0;
                       end 
                      
                  10'sd150/*150:xpc10*/:  begin 
                       xpc10 <= 10'sd151/*151:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'shda] <= 8'h0;
                       A_8_US_CC_SCALbx14_ARA0[64'shd9] <= 8'h0;
                       end 
                      
                  10'sd151/*151:xpc10*/:  begin 
                       xpc10 <= 10'sd152/*152:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'shdc] <= 8'h0;
                       A_8_US_CC_SCALbx14_ARA0[64'shdb] <= 8'h0;
                       end 
                      
                  10'sd152/*152:xpc10*/:  begin 
                       xpc10 <= 10'sd153/*153:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'shde] <= 8'h0;
                       A_8_US_CC_SCALbx14_ARA0[64'shdd] <= 8'h0;
                       end 
                      
                  10'sd153/*153:xpc10*/:  begin 
                       xpc10 <= 10'sd154/*154:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'she0] <= 8'h0;
                       A_8_US_CC_SCALbx14_ARA0[64'shdf] <= 8'h0;
                       end 
                      
                  10'sd154/*154:xpc10*/:  begin 
                       xpc10 <= 10'sd155/*155:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'she2] <= 8'h0;
                       A_8_US_CC_SCALbx14_ARA0[64'she1] <= 8'h0;
                       end 
                      
                  10'sd155/*155:xpc10*/:  begin 
                       xpc10 <= 10'sd156/*156:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'she4] <= 8'h0;
                       A_8_US_CC_SCALbx14_ARA0[64'she3] <= 8'h0;
                       end 
                      
                  10'sd156/*156:xpc10*/:  begin 
                       xpc10 <= 10'sd157/*157:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'she6] <= 8'h0;
                       A_8_US_CC_SCALbx14_ARA0[64'she5] <= 8'h0;
                       end 
                      
                  10'sd157/*157:xpc10*/:  begin 
                       xpc10 <= 10'sd158/*158:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'she8] <= 8'h0;
                       A_8_US_CC_SCALbx14_ARA0[64'she7] <= 8'h0;
                       end 
                      
                  10'sd158/*158:xpc10*/:  begin 
                       xpc10 <= 10'sd159/*159:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'shea] <= 8'h0;
                       A_8_US_CC_SCALbx14_ARA0[64'she9] <= 8'h0;
                       end 
                      
                  10'sd159/*159:xpc10*/:  begin 
                       xpc10 <= 10'sd160/*160:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'shec] <= 8'h0;
                       A_8_US_CC_SCALbx14_ARA0[64'sheb] <= 8'h0;
                       end 
                      
                  10'sd160/*160:xpc10*/:  begin 
                       xpc10 <= 10'sd161/*161:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'shee] <= 8'h0;
                       A_8_US_CC_SCALbx14_ARA0[64'shed] <= 8'h0;
                       end 
                      
                  10'sd161/*161:xpc10*/:  begin 
                       xpc10 <= 10'sd162/*162:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'shf0] <= 8'h0;
                       A_8_US_CC_SCALbx14_ARA0[64'shef] <= 8'h0;
                       end 
                      
                  10'sd162/*162:xpc10*/:  begin 
                       xpc10 <= 10'sd163/*163:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'shf2] <= 8'h0;
                       A_8_US_CC_SCALbx14_ARA0[64'shf1] <= 8'h0;
                       end 
                      
                  10'sd163/*163:xpc10*/:  begin 
                       xpc10 <= 10'sd164/*164:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'shf4] <= 8'h0;
                       A_8_US_CC_SCALbx14_ARA0[64'shf3] <= 8'h0;
                       end 
                      
                  10'sd164/*164:xpc10*/:  begin 
                       xpc10 <= 10'sd165/*165:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'shf6] <= 8'h0;
                       A_8_US_CC_SCALbx14_ARA0[64'shf5] <= 8'h0;
                       end 
                      
                  10'sd165/*165:xpc10*/:  begin 
                       xpc10 <= 10'sd166/*166:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'shf8] <= 8'h0;
                       A_8_US_CC_SCALbx14_ARA0[64'shf7] <= 8'h0;
                       end 
                      
                  10'sd166/*166:xpc10*/:  begin 
                       xpc10 <= 10'sd167/*167:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'shfa] <= 8'h0;
                       A_8_US_CC_SCALbx14_ARA0[64'shf9] <= 8'h0;
                       end 
                      
                  10'sd167/*167:xpc10*/:  begin 
                       xpc10 <= 10'sd168/*168:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'shfc] <= 8'h0;
                       A_8_US_CC_SCALbx14_ARA0[64'shfb] <= 8'h0;
                       end 
                      
                  10'sd168/*168:xpc10*/:  begin 
                       xpc10 <= 10'sd169/*169:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'shfe] <= 8'h0;
                       A_8_US_CC_SCALbx14_ARA0[64'shfd] <= 8'h0;
                       end 
                      
                  10'sd169/*169:xpc10*/:  begin 
                       xpc10 <= 10'sd170/*170:xpc10*/;
                       A_8_US_CC_SCALbx14_ARA0[64'shff] <= 8'h0;
                       end 
                      
                  10'sd171/*171:xpc10*/:  xpc10 <= 10'sd172/*172:xpc10*/;

                  10'sd172/*172:xpc10*/:  begin 
                       xpc10 <= 10'sd173/*173:xpc10*/;
                       Tdbm0_3_V_1 <= 32'sd0;
                       Tdbm0_3_V_0 <= 32'sd0;
                       end 
                      
                  10'sd174/*174:xpc10*/:  begin 
                       xpc10 <= 10'sd175/*175:xpc10*/;
                       Tdsi3_5_V_0 <= $unsigned(A_64_US_CC_SCALbx12_ARB0[Tdbm0_3_V_1]);
                       end 
                      
                  10'sd175/*175:xpc10*/:  begin 
                       xpc10 <= 10'sd176/*176:xpc10*/;
                       Tdsi3_5_V_1 <= $unsigned(A_64_US_CC_SCALbx12_ARB0[Tdbm0_3_V_1]);
                       end 
                      
                  10'sd176/*176:xpc10*/:  begin 
                       xpc10 <= 10'sd177/*177:xpc10*/;
                       Tsfl0_9_V_8 <= 64'h0;
                       Tdsi3_5_V_2 <= 32'sd1;
                       end 
                      
                  10'sd177/*177:xpc10*/:  begin 
                       xpc10 <= 10'sd178/*178:xpc10*/;
                       Tsfl0_9_V_6 <= 64'shf_ffff_ffff_ffff&A_64_US_CC_SCALbx12_ARB0[Tdbm0_3_V_1];
                       Tsfl0_9_V_9 <= 64'h0;
                       end 
                      
                  10'sd178/*178:xpc10*/:  begin 
                       xpc10 <= 10'sd179/*179:xpc10*/;
                       Tsfl0_9_V_3 <= rtl_signed_bitextract9(64'sh7ff&(A_64_US_CC_SCALbx12_ARB0[Tdbm0_3_V_1]>>32'sd52));
                       end 
                      
                  10'sd180/*180:xpc10*/:  begin 
                       xpc10 <= 10'sd181/*181:xpc10*/;
                       Tsfl0_9_V_7 <= 64'shf_ffff_ffff_ffff&A_64_US_CC_SCALbx12_ARB0[Tdbm0_3_V_1];
                       end 
                      
                  10'sd181/*181:xpc10*/:  begin 
                       xpc10 <= 10'sd182/*182:xpc10*/;
                       Tsfl0_9_V_4 <= rtl_signed_bitextract9(64'sh7ff&(A_64_US_CC_SCALbx12_ARB0[Tdbm0_3_V_1]>>32'sd52));
                       end 
                      
                  10'sd183/*183:xpc10*/:  begin 
                       xpc10 <= 10'sd184/*184:xpc10*/;
                       Tsfl0_9_V_2 <= rtl_unsigned_bitextract8(Tsfl0_9_V_0^Tsfl0_9_V_1);
                       end 
                      
                  10'sd185/*185:xpc10*/:  begin 
                       xpc10 <= 10'sd186/*186:xpc10*/;
                       Tspr4_3_V_1 <= $unsigned(A_64_US_CC_SCALbx12_ARB0[Tdbm0_3_V_1]);
                       end 
                      
                  10'sd187/*187:xpc10*/:  begin 
                       xpc10 <= 10'sd188/*188:xpc10*/;
                       Tspr4_3_V_3 <= (-64'sh20_0000_0000_0000<$signed((Tspr4_3_V_1<<32'sd1)));
                       Tspr4_3_V_2 <= rtl_unsigned_bitextract5(Tsf0SPILL10_256);
                       end 
                      
                  10'sd189/*189:xpc10*/:  begin 
                       xpc10 <= 10'sd190/*190:xpc10*/;
                       Tspr4_3_V_0 <= 64'sh8_0000_0000_0000|Tspr4_3_V_0;
                       Tspr4_3_V_4 <= rtl_unsigned_bitextract5(Tsf0SPILL12_256);
                       end 
                      
                  10'sd190/*190:xpc10*/:  begin 
                       xpc10 <= 10'sd191/*191:xpc10*/;
                       Tspr4_3_V_1 <= 64'sh8_0000_0000_0000|Tspr4_3_V_1;
                       end 
                      
                  10'sd193/*193:xpc10*/:  begin 
                       xpc10 <= 10'sd194/*194:xpc10*/;
                       Tsfl0_10_V_0 <= -64'sh_8000_0000_0000_0000&~Tsf0_SPILL_256|64'sh_7fff_ffff_ffff_ffff&Tsf0_SPILL_256;
                       end 
                      
                  10'sd194/*194:xpc10*/:  begin 
                       xpc10 <= 10'sd195/*195:xpc10*/;
                       dfsin_gloops <= 32'sd1+dfsin_gloops;
                       Tdsi3_5_V_3 <= Tsfl0_10_V_0;
                       end 
                      
                  10'sd195/*195:xpc10*/:  begin 
                       xpc10 <= 10'sd196/*196:xpc10*/;
                       Tsfl1_7_V_9 <= 64'h0;
                       Tsfl1_7_V_8 <= 64'h0;
                       end 
                      
                  10'sd196/*196:xpc10*/:  begin 
                       xpc10 <= 10'sd197/*197:xpc10*/;
                       Tsfl1_7_V_6 <= 64'shf_ffff_ffff_ffff&Tdsi3_5_V_1;
                       end 
                      
                  10'sd197/*197:xpc10*/:  begin 
                       xpc10 <= 10'sd198/*198:xpc10*/;
                       Tsfl1_7_V_3 <= rtl_signed_bitextract9(64'sh7ff&(Tdsi3_5_V_1>>32'sd52));
                       end 
                      
                  10'sd199/*199:xpc10*/:  begin 
                       xpc10 <= 10'sd200/*200:xpc10*/;
                       Tsfl1_7_V_7 <= 64'shf_ffff_ffff_ffff&Tdsi3_5_V_3;
                       end 
                      
                  10'sd200/*200:xpc10*/:  begin 
                       xpc10 <= 10'sd201/*201:xpc10*/;
                       Tsfl1_7_V_4 <= rtl_signed_bitextract9(64'sh7ff&(Tdsi3_5_V_3>>32'sd52));
                       end 
                      
                  10'sd201/*201:xpc10*/: if ((64'sh0<(Tdsi3_5_V_3>>32'sd63)))  begin 
                           xpc10 <= 10'sd202/*202:xpc10*/;
                           Tsfl1_7_V_1 <= 1'h1;
                           end 
                           else  begin 
                           xpc10 <= 10'sd202/*202:xpc10*/;
                           Tsfl1_7_V_1 <= 1'h0;
                           end 
                          
                  10'sd202/*202:xpc10*/:  begin 
                       xpc10 <= 10'sd203/*203:xpc10*/;
                       Tsfl1_7_V_2 <= rtl_unsigned_bitextract8(Tsfl1_7_V_0^Tsfl1_7_V_1);
                       end 
                      
                  10'sd205/*205:xpc10*/:  begin 
                       xpc10 <= 10'sd206/*206:xpc10*/;
                       Tspr4_3_V_3 <= (-64'sh20_0000_0000_0000<$signed((Tspr4_3_V_1<<32'sd1)));
                       Tspr4_3_V_2 <= rtl_unsigned_bitextract5(Tsf0SPILL10_256);
                       end 
                      
                  10'sd207/*207:xpc10*/:  begin 
                       xpc10 <= 10'sd208/*208:xpc10*/;
                       Tspr4_3_V_0 <= 64'sh8_0000_0000_0000|Tspr4_3_V_0;
                       Tspr4_3_V_4 <= rtl_unsigned_bitextract5(Tsf0SPILL12_256);
                       end 
                      
                  10'sd208/*208:xpc10*/:  begin 
                       xpc10 <= 10'sd209/*209:xpc10*/;
                       Tspr4_3_V_1 <= 64'sh8_0000_0000_0000|Tspr4_3_V_1;
                       end 
                      
                  10'sd212/*212:xpc10*/:  begin 
                       xpc10 <= 10'sd213/*213:xpc10*/;
                       Tsfl1_18_V_3 <= rtl_signed_bitextract9(64'sh7ff&(Tsf1_SPILL_256>>32'sd52));
                       end 
                      
                  10'sd213/*213:xpc10*/: if ((64'sh0<(Tsf1_SPILL_256>>32'sd63)))  begin 
                           xpc10 <= 10'sd214/*214:xpc10*/;
                           Tsfl1_18_V_0 <= 1'h1;
                           end 
                           else  begin 
                           xpc10 <= 10'sd214/*214:xpc10*/;
                           Tsfl1_18_V_0 <= 1'h0;
                           end 
                          
                  10'sd214/*214:xpc10*/:  begin 
                       xpc10 <= 10'sd215/*215:xpc10*/;
                       Tsfl1_18_V_7 <= 64'shf_ffff_ffff_ffff&Tsi1_SPILL_256;
                       end 
                      
                  10'sd215/*215:xpc10*/:  begin 
                       xpc10 <= 10'sd216/*216:xpc10*/;
                       Tsfl1_18_V_4 <= rtl_signed_bitextract9(64'sh7ff&(Tsi1_SPILL_256>>32'sd52));
                       end 
                      
                  10'sd216/*216:xpc10*/: if ((64'sh0<(Tsi1_SPILL_256>>32'sd63)))  begin 
                           xpc10 <= 10'sd217/*217:xpc10*/;
                           Tsfl1_18_V_1 <= 1'h1;
                           end 
                           else  begin 
                           xpc10 <= 10'sd217/*217:xpc10*/;
                           Tsfl1_18_V_1 <= 1'h0;
                           end 
                          
                  10'sd217/*217:xpc10*/:  begin 
                       xpc10 <= 10'sd218/*218:xpc10*/;
                       Tsfl1_18_V_2 <= rtl_unsigned_bitextract8(Tsfl1_18_V_0^Tsfl1_18_V_1);
                       end 
                      
                  10'sd220/*220:xpc10*/:  begin 
                       xpc10 <= 10'sd221/*221:xpc10*/;
                       Tspr2_2_V_3 <= (-64'sh20_0000_0000_0000<$signed((Tspr2_2_V_1<<32'sd1)));
                       Tspr2_2_V_2 <= rtl_unsigned_bitextract5(Tsf0SPILL10_256);
                       end 
                      
                  10'sd222/*222:xpc10*/:  begin 
                       xpc10 <= 10'sd223/*223:xpc10*/;
                       Tspr2_2_V_0 <= 64'sh8_0000_0000_0000|Tspr2_2_V_0;
                       Tspr2_2_V_4 <= rtl_unsigned_bitextract5(Tsf0SPILL12_256);
                       end 
                      
                  10'sd223/*223:xpc10*/:  begin 
                       xpc10 <= 10'sd224/*224:xpc10*/;
                       Tspr2_2_V_1 <= 64'sh8_0000_0000_0000|Tspr2_2_V_1;
                       end 
                      
                  10'sd229/*229:xpc10*/:  begin 
                       xpc10 <= 10'sd230/*230:xpc10*/;
                       Tsad1_3_V_0 <= rtl_signed_bitextract9(64'sh7ff&(Tdsi3_5_V_0>>32'sd52));
                       end 
                      
                  10'sd230/*230:xpc10*/:  begin 
                       xpc10 <= 10'sd231/*231:xpc10*/;
                       Tsad1_3_V_4 <= 64'shf_ffff_ffff_ffff&Tdsi3_5_V_1;
                       end 
                      
                  10'sd231/*231:xpc10*/:  begin 
                       xpc10 <= 10'sd232/*232:xpc10*/;
                       Tsad1_3_V_1 <= rtl_signed_bitextract9(64'sh7ff&(Tdsi3_5_V_1>>32'sd52));
                       end 
                      
                  10'sd232/*232:xpc10*/:  begin 
                       xpc10 <= 10'sd233/*233:xpc10*/;
                       Tsad1_3_V_6 <= rtl_sign_extend2(Tsad1_3_V_0)+(0-Tsad1_3_V_1);
                       end 
                      
                  10'sd233/*233:xpc10*/:  begin 
                       xpc10 <= 10'sd234/*234:xpc10*/;
                       Tsad1_3_V_3 <= (Tsad1_3_V_3<<32'sd9);
                       end 
                      
                  10'sd234/*234:xpc10*/:  begin 
                       xpc10 <= 10'sd235/*235:xpc10*/;
                       Tsad1_3_V_4 <= (Tsad1_3_V_4<<32'sd9);
                       end 
                      
                  10'sd237/*237:xpc10*/:  begin 
                       xpc10 <= 10'sd238/*238:xpc10*/;
                       Tspr3_2_V_3 <= (-64'sh20_0000_0000_0000<$signed((Tspr3_2_V_1<<32'sd1)));
                       Tspr3_2_V_2 <= rtl_unsigned_bitextract5(Tsf0SPILL10_256);
                       end 
                      
                  10'sd239/*239:xpc10*/:  begin 
                       xpc10 <= 10'sd240/*240:xpc10*/;
                       Tspr3_2_V_0 <= 64'sh8_0000_0000_0000|Tspr3_2_V_0;
                       Tspr3_2_V_4 <= rtl_unsigned_bitextract5(Tsf0SPILL12_256);
                       end 
                      
                  10'sd240/*240:xpc10*/:  begin 
                       xpc10 <= 10'sd241/*241:xpc10*/;
                       Tspr3_2_V_1 <= 64'sh8_0000_0000_0000|Tspr3_2_V_1;
                       end 
                      
                  10'sd243/*243:xpc10*/:  begin 
                       xpc10 <= 10'sd244/*244:xpc10*/;
                       Tdsi3_5_V_0 <= Tsa1_SPILL_256;
                       Tsf1SPILL12_256 <= Tsa1_SPILL_256;
                       end 
                      
                  10'sd244/*244:xpc10*/:  begin 
                       xpc10 <= 10'sd245/*245:xpc10*/;
                       Tdsi3_5_V_2 <= 32'sd1+Tdsi3_5_V_2;
                       end 
                      
                  10'sd246/*246:xpc10*/:  begin 
                       xpc10 <= 10'sd247/*247:xpc10*/;
                       Tdbm0_3_V_2 <= Tdsi3_5_V_0;
                       Tsf0SPILL14_256 <= 32'sd0;
                       end 
                      
                  10'sd247/*247:xpc10*/:  begin 
                       xpc10 <= 10'sd248/*248:xpc10*/;
                       Tdb0_SPILL_259 <= Tdbm0_3_V_0;
                       fastspilldup76 <= Tdbm0_3_V_0;
                       end 
                      
                  10'sd249/*249:xpc10*/:  begin 
                       xpc10 <= 10'sd250/*250:xpc10*/;
                       Tdbm0_3_V_0 <= Tdb0_SPILL_256+Tdb0_SPILL_258;
                       end 
                      
                  10'sd250/*250:xpc10*/:  xpc10 <= 10'sd251/*251:xpc10*/;

                  10'sd252/*252:xpc10*/:  begin 
                       xpc10 <= 10'sd253/*253:xpc10*/;
                       Tdbm0_3_V_1 <= 32'sd1+Tdbm0_3_V_1;
                       end 
                      
                  10'sd257/*257:xpc10*/:  begin 
                       xpc10 <= 10'sd250/*250:xpc10*/;
                       Tdbm0_3_V_0 <= Tdb0_SPILL_259+Tdb0_SPILL_258;
                       end 
                      
                  10'sd264/*264:xpc10*/:  begin 
                       xpc10 <= 10'sd240/*240:xpc10*/;
                       Tspr3_2_V_0 <= 64'sh8_0000_0000_0000|Tspr3_2_V_0;
                       end 
                      
                  10'sd265/*265:xpc10*/:  begin 
                       xpc10 <= 10'sd238/*238:xpc10*/;
                       Tspr3_2_V_3 <= (-64'sh20_0000_0000_0000<$signed((Tspr3_2_V_1<<32'sd1)));
                       end 
                      
                  10'sd266/*266:xpc10*/:  begin 
                       xpc10 <= 10'sd245/*245:xpc10*/;
                       Tdsi3_5_V_2 <= 32'sd1+Tdsi3_5_V_2;
                       Tdsi3_5_V_0 <= Tsf1SPILL12_256;
                       end 
                      
                  10'sd268/*268:xpc10*/:  begin 
                       xpc10 <= 10'sd269/*269:xpc10*/;
                       Tsad1_3_V_3 <= 64'sh_2000_0000_0000_0000|Tsad1_3_V_3;
                       Tsad1_3_V_2 <= rtl_signed_bitextract0(Tsad1_3_V_0);
                       end 
                      
                  10'sd269/*269:xpc10*/:  begin 
                       xpc10 <= 10'sd270/*270:xpc10*/;
                       Tsad1_3_V_5 <= (Tsad1_3_V_3+Tsad1_3_V_4<<32'sd1);
                       end 
                      
                  10'sd270/*270:xpc10*/:  begin 
                       xpc10 <= 10'sd271/*271:xpc10*/;
                       Tsad1_3_V_2 <= rtl_signed_bitextract0(-16'sd1+Tsad1_3_V_2);
                       end 
                      
                  10'sd272/*272:xpc10*/:  begin 
                       xpc10 <= 10'sd273/*273:xpc10*/;
                       Tsad1_3_V_2 <= rtl_signed_bitextract0(16'sd1+Tsad1_3_V_2);
                       end 
                      
                  10'sd273/*273:xpc10*/:  begin 
                       xpc10 <= 10'sd274/*274:xpc10*/;
                       Tsro28_4_V_1 <= Tsad1_3_V_5;
                       Tsro28_4_V_0 <= rtl_signed_bitextract0(Tsad1_3_V_2);
                       end 
                      
                  10'sd275/*275:xpc10*/:  begin 
                       xpc10 <= 10'sd276/*276:xpc10*/;
                       Tsro28_4_V_6 <= rtl_signed_bitextract9(64'sh3ff&Tsro28_4_V_1);
                       Tsro28_4_V_5 <= 16'sh200;
                       end 
                      
                  10'sd278/*278:xpc10*/:  begin 
                       xpc10 <= 10'sd279/*279:xpc10*/;
                       Tsr28_SPILL_256 <= fastspilldup64;
                       Tsr28_SPILL_260 <= fastspilldup64;
                       end 
                      
                  10'sd280/*280:xpc10*/:  begin 
                       xpc10 <= 10'sd281/*281:xpc10*/;
                       Tsr28_SPILL_259 <= Tsr28_SPILL_257+(0-Tsr28_SPILL_258);
                       end 
                      
                  10'sd281/*281:xpc10*/:  begin 
                       xpc10 <= 10'sd266/*266:xpc10*/;
                       Tsf1SPILL12_256 <= Tsr28_SPILL_259;
                       Tsa1_SPILL_256 <= Tsr28_SPILL_259;
                       end 
                      
                  10'sd282/*282:xpc10*/:  begin 
                       xpc10 <= 10'sd281/*281:xpc10*/;
                       Tsr28_SPILL_259 <= Tsr28_SPILL_257+(0-Tsr28_SPILL_258);
                       end 
                      
                  10'sd283/*283:xpc10*/:  begin 
                       xpc10 <= 10'sd284/*284:xpc10*/;
                       Tsro28_4_V_0 <= 16'sh0;
                       Tsro28_4_V_1 <= Tssh18_7_V_0;
                       end 
                      
                  10'sd284/*284:xpc10*/:  begin 
                       xpc10 <= 10'sd285/*285:xpc10*/;
                       Tsro28_4_V_6 <= rtl_signed_bitextract9(64'sh3ff&Tsro28_4_V_1);
                       end 
                      
                  10'sd287/*287:xpc10*/:  begin 
                       xpc10 <= 10'sd288/*288:xpc10*/;
                       Tsro28_4_V_1 <= (Tsro28_4_V_1+rtl_sign_extend4(Tsro28_4_V_5)>>32'sd10);
                       end 
                      
                  10'sd290/*290:xpc10*/:  begin 
                       xpc10 <= 10'sd291/*291:xpc10*/;
                       Tsr28_SPILL_259 <= Tsro28_4_V_1+(Tsp27_SPILL_256<<32'sd63)+(rtl_sign_extend4(Tsro28_4_V_0)<<32'sd52);
                       end 
                      
                  10'sd291/*291:xpc10*/:  begin 
                       xpc10 <= 10'sd266/*266:xpc10*/;
                       Tsf1SPILL12_256 <= Tsr28_SPILL_259;
                       Tsa1_SPILL_256 <= Tsr28_SPILL_259;
                       end 
                      
                  10'sd292/*292:xpc10*/:  begin 
                       xpc10 <= 10'sd291/*291:xpc10*/;
                       Tsr28_SPILL_259 <= Tsro28_4_V_1+(Tsp27_SPILL_256<<32'sd63)+(rtl_sign_extend4(Tsro28_4_V_0)<<32'sd52);
                       end 
                      
                  10'sd293/*293:xpc10*/:  begin 
                       xpc10 <= 10'sd294/*294:xpc10*/;
                       Tss18_SPILL_256 <= fastspilldup66;
                       Tss18_SPILL_259 <= fastspilldup66;
                       end 
                      
                  10'sd295/*295:xpc10*/:  begin 
                       xpc10 <= 10'sd296/*296:xpc10*/;
                       Tssh18_7_V_0 <= Tss18_SPILL_258|Tss18_SPILL_257;
                       end 
                      
                  10'sd296/*296:xpc10*/:  begin 
                       xpc10 <= 10'sd284/*284:xpc10*/;
                       Tsro28_4_V_0 <= 16'sh0;
                       Tsro28_4_V_1 <= Tssh18_7_V_0;
                       end 
                      
                  10'sd297/*297:xpc10*/:  begin 
                       xpc10 <= 10'sd296/*296:xpc10*/;
                       Tssh18_7_V_0 <= Tss18_SPILL_258|Tss18_SPILL_257;
                       end 
                      
                  10'sd298/*298:xpc10*/:  begin 
                       xpc10 <= 10'sd299/*299:xpc10*/;
                       Tsro28_4_V_1 <= Tss18_SPILL_260;
                       Tssh18_7_V_0 <= Tss18_SPILL_260;
                       end 
                      
                  10'sd299/*299:xpc10*/:  begin 
                       xpc10 <= 10'sd285/*285:xpc10*/;
                       Tsro28_4_V_6 <= rtl_signed_bitextract9(64'sh3ff&Tsro28_4_V_1);
                       Tsro28_4_V_0 <= 16'sh0;
                       end 
                      
                  10'sd300/*300:xpc10*/:  begin 
                       xpc10 <= 10'sd299/*299:xpc10*/;
                       Tsro28_4_V_1 <= Tss18_SPILL_260;
                       Tssh18_7_V_0 <= Tss18_SPILL_260;
                       end 
                      
                  10'sd301/*301:xpc10*/:  begin 
                       xpc10 <= 10'sd302/*302:xpc10*/;
                       Tss8_SPILL_256 <= fastspilldup60;
                       Tss8_SPILL_259 <= fastspilldup60;
                       end 
                      
                  10'sd303/*303:xpc10*/:  begin 
                       xpc10 <= 10'sd304/*304:xpc10*/;
                       Tssh8_5_V_0 <= Tss8_SPILL_258|Tss8_SPILL_257;
                       end 
                      
                  10'sd304/*304:xpc10*/:  begin 
                       xpc10 <= 10'sd305/*305:xpc10*/;
                       Tsad1_3_V_2 <= rtl_signed_bitextract0(Tsad1_3_V_0);
                       Tsad1_3_V_4 <= Tssh8_5_V_0;
                       end 
                      
                  10'sd305/*305:xpc10*/:  begin 
                       xpc10 <= 10'sd269/*269:xpc10*/;
                       Tsad1_3_V_3 <= 64'sh_2000_0000_0000_0000|Tsad1_3_V_3;
                       end 
                      
                  10'sd306/*306:xpc10*/:  begin 
                       xpc10 <= 10'sd304/*304:xpc10*/;
                       Tssh8_5_V_0 <= Tss8_SPILL_258|Tss8_SPILL_257;
                       end 
                      
                  10'sd307/*307:xpc10*/:  begin 
                       xpc10 <= 10'sd305/*305:xpc10*/;
                       Tsad1_3_V_2 <= rtl_signed_bitextract0(Tsad1_3_V_0);
                       Tsad1_3_V_4 <= Tssh8_5_V_0;
                       end 
                      
                  10'sd310/*310:xpc10*/:  begin 
                       xpc10 <= 10'sd311/*311:xpc10*/;
                       Tspr12_2_V_3 <= (-64'sh20_0000_0000_0000<$signed((Tspr12_2_V_1<<32'sd1)));
                       Tspr12_2_V_2 <= rtl_unsigned_bitextract5(Tsf0SPILL10_256);
                       end 
                      
                  10'sd312/*312:xpc10*/:  begin 
                       xpc10 <= 10'sd313/*313:xpc10*/;
                       Tspr12_2_V_0 <= 64'sh8_0000_0000_0000|Tspr12_2_V_0;
                       Tspr12_2_V_4 <= rtl_unsigned_bitextract5(Tsf0SPILL12_256);
                       end 
                      
                  10'sd313/*313:xpc10*/:  begin 
                       xpc10 <= 10'sd314/*314:xpc10*/;
                       Tspr12_2_V_1 <= 64'sh8_0000_0000_0000|Tspr12_2_V_1;
                       end 
                      
                  10'sd316/*316:xpc10*/:  begin 
                       xpc10 <= 10'sd244/*244:xpc10*/;
                       Tdsi3_5_V_0 <= Tsa1_SPILL_256;
                       Tsf1SPILL12_256 <= Tsa1_SPILL_256;
                       end 
                      
                  10'sd317/*317:xpc10*/:  begin 
                       xpc10 <= 10'sd313/*313:xpc10*/;
                       Tspr12_2_V_0 <= 64'sh8_0000_0000_0000|Tspr12_2_V_0;
                       end 
                      
                  10'sd318/*318:xpc10*/:  begin 
                       xpc10 <= 10'sd311/*311:xpc10*/;
                       Tspr12_2_V_3 <= (-64'sh20_0000_0000_0000<$signed((Tspr12_2_V_1<<32'sd1)));
                       end 
                      
                  10'sd319/*319:xpc10*/:  begin 
                       xpc10 <= 10'sd244/*244:xpc10*/;
                       Tdsi3_5_V_0 <= Tsa1_SPILL_256;
                       Tsf1SPILL12_256 <= Tsa1_SPILL_256;
                       end 
                      
                  10'sd321/*321:xpc10*/:  begin 
                       xpc10 <= 10'sd269/*269:xpc10*/;
                       Tsad1_3_V_3 <= 64'sh_2000_0000_0000_0000|Tsad1_3_V_3;
                       Tsad1_3_V_2 <= rtl_signed_bitextract0(Tsad1_3_V_1);
                       end 
                      
                  10'sd322/*322:xpc10*/:  begin 
                       xpc10 <= 10'sd323/*323:xpc10*/;
                       Tss17_SPILL_256 <= fastspilldup62;
                       Tss17_SPILL_259 <= fastspilldup62;
                       end 
                      
                  10'sd324/*324:xpc10*/:  begin 
                       xpc10 <= 10'sd325/*325:xpc10*/;
                       Tssh17_6_V_0 <= Tss17_SPILL_258|Tss17_SPILL_257;
                       end 
                      
                  10'sd325/*325:xpc10*/:  begin 
                       xpc10 <= 10'sd326/*326:xpc10*/;
                       Tsad1_3_V_2 <= rtl_signed_bitextract0(Tsad1_3_V_1);
                       Tsad1_3_V_3 <= Tssh17_6_V_0;
                       end 
                      
                  10'sd326/*326:xpc10*/:  begin 
                       xpc10 <= 10'sd269/*269:xpc10*/;
                       Tsad1_3_V_3 <= 64'sh_2000_0000_0000_0000|Tsad1_3_V_3;
                       end 
                      
                  10'sd327/*327:xpc10*/:  begin 
                       xpc10 <= 10'sd325/*325:xpc10*/;
                       Tssh17_6_V_0 <= Tss17_SPILL_258|Tss17_SPILL_257;
                       end 
                      
                  10'sd328/*328:xpc10*/:  begin 
                       xpc10 <= 10'sd326/*326:xpc10*/;
                       Tsad1_3_V_2 <= rtl_signed_bitextract0(Tsad1_3_V_1);
                       Tsad1_3_V_3 <= Tssh17_6_V_0;
                       end 
                      
                  10'sd331/*331:xpc10*/:  begin 
                       xpc10 <= 10'sd332/*332:xpc10*/;
                       Tspr21_3_V_3 <= (-64'sh20_0000_0000_0000<$signed((Tspr21_3_V_1<<32'sd1)));
                       Tspr21_3_V_2 <= rtl_unsigned_bitextract5(Tsf0SPILL10_256);
                       end 
                      
                  10'sd333/*333:xpc10*/:  begin 
                       xpc10 <= 10'sd334/*334:xpc10*/;
                       Tspr21_3_V_0 <= 64'sh8_0000_0000_0000|Tspr21_3_V_0;
                       Tspr21_3_V_4 <= rtl_unsigned_bitextract5(Tsf0SPILL12_256);
                       end 
                      
                  10'sd334/*334:xpc10*/:  begin 
                       xpc10 <= 10'sd335/*335:xpc10*/;
                       Tspr21_3_V_1 <= 64'sh8_0000_0000_0000|Tspr21_3_V_1;
                       end 
                      
                  10'sd337/*337:xpc10*/:  begin 
                       xpc10 <= 10'sd244/*244:xpc10*/;
                       Tdsi3_5_V_0 <= Tsa1_SPILL_256;
                       Tsf1SPILL12_256 <= Tsa1_SPILL_256;
                       end 
                      
                  10'sd338/*338:xpc10*/:  begin 
                       xpc10 <= 10'sd334/*334:xpc10*/;
                       Tspr21_3_V_0 <= 64'sh8_0000_0000_0000|Tspr21_3_V_0;
                       end 
                      
                  10'sd339/*339:xpc10*/:  begin 
                       xpc10 <= 10'sd332/*332:xpc10*/;
                       Tspr21_3_V_3 <= (-64'sh20_0000_0000_0000<$signed((Tspr21_3_V_1<<32'sd1)));
                       end 
                      
                  10'sd340/*340:xpc10*/:  begin 
                       xpc10 <= 10'sd244/*244:xpc10*/;
                       Tdsi3_5_V_0 <= Tsa1_SPILL_256;
                       Tsf1SPILL12_256 <= Tsa1_SPILL_256;
                       end 
                      
                  10'sd341/*341:xpc10*/:  begin 
                       xpc10 <= 10'sd342/*342:xpc10*/;
                       Tsro28_4_V_0 <= rtl_signed_bitextract0(Tsad1_3_V_0);
                       Tsad1_3_V_2 <= rtl_signed_bitextract0(Tsad1_3_V_0);
                       end 
                      
                  10'sd342/*342:xpc10*/:  begin 
                       xpc10 <= 10'sd343/*343:xpc10*/;
                       Tsro28_4_V_1 <= Tsad1_3_V_5;
                       end 
                      
                  10'sd343/*343:xpc10*/:  begin 
                       xpc10 <= 10'sd344/*344:xpc10*/;
                       Tsro28_4_V_5 <= 16'sh200;
                       end 
                      
                  10'sd344/*344:xpc10*/:  begin 
                       xpc10 <= 10'sd276/*276:xpc10*/;
                       Tsro28_4_V_6 <= rtl_signed_bitextract9(64'sh3ff&Tsro28_4_V_1);
                       end 
                      
                  10'sd345/*345:xpc10*/:  begin 
                       xpc10 <= 10'sd346/*346:xpc10*/;
                       Tssu2_4_V_4 <= 64'shf_ffff_ffff_ffff&Tdsi3_5_V_0;
                       end 
                      
                  10'sd346/*346:xpc10*/:  begin 
                       xpc10 <= 10'sd347/*347:xpc10*/;
                       Tssu2_4_V_1 <= rtl_signed_bitextract9(64'sh7ff&(Tdsi3_5_V_0>>32'sd52));
                       end 
                      
                  10'sd347/*347:xpc10*/:  begin 
                       xpc10 <= 10'sd348/*348:xpc10*/;
                       Tssu2_4_V_5 <= 64'shf_ffff_ffff_ffff&Tdsi3_5_V_1;
                       end 
                      
                  10'sd348/*348:xpc10*/:  begin 
                       xpc10 <= 10'sd349/*349:xpc10*/;
                       Tssu2_4_V_2 <= rtl_signed_bitextract9(64'sh7ff&(Tdsi3_5_V_1>>32'sd52));
                       end 
                      
                  10'sd349/*349:xpc10*/:  begin 
                       xpc10 <= 10'sd350/*350:xpc10*/;
                       Tssu2_4_V_7 <= rtl_sign_extend2(Tssu2_4_V_1)+(0-Tssu2_4_V_2);
                       end 
                      
                  10'sd350/*350:xpc10*/:  begin 
                       xpc10 <= 10'sd351/*351:xpc10*/;
                       Tssu2_4_V_4 <= (Tssu2_4_V_4<<32'sd10);
                       end 
                      
                  10'sd351/*351:xpc10*/:  begin 
                       xpc10 <= 10'sd352/*352:xpc10*/;
                       Tssu2_4_V_5 <= (Tssu2_4_V_5<<32'sd10);
                       end 
                      
                  10'sd354/*354:xpc10*/:  begin 
                       xpc10 <= 10'sd355/*355:xpc10*/;
                       Tspr27_2_V_3 <= (-64'sh20_0000_0000_0000<$signed((Tspr27_2_V_1<<32'sd1)));
                       Tspr27_2_V_2 <= rtl_unsigned_bitextract5(Tsf0SPILL10_256);
                       end 
                      
                  10'sd356/*356:xpc10*/:  begin 
                       xpc10 <= 10'sd357/*357:xpc10*/;
                       Tspr27_2_V_0 <= 64'sh8_0000_0000_0000|Tspr27_2_V_0;
                       Tspr27_2_V_4 <= rtl_unsigned_bitextract5(Tsf0SPILL12_256);
                       end 
                      
                  10'sd357/*357:xpc10*/:  begin 
                       xpc10 <= 10'sd358/*358:xpc10*/;
                       Tspr27_2_V_1 <= 64'sh8_0000_0000_0000|Tspr27_2_V_1;
                       end 
                      
                  10'sd360/*360:xpc10*/:  begin 
                       xpc10 <= 10'sd244/*244:xpc10*/;
                       Tdsi3_5_V_0 <= Tss2_SPILL_256;
                       Tsf1SPILL12_256 <= Tss2_SPILL_256;
                       end 
                      
                  10'sd361/*361:xpc10*/:  begin 
                       xpc10 <= 10'sd357/*357:xpc10*/;
                       Tspr27_2_V_0 <= 64'sh8_0000_0000_0000|Tspr27_2_V_0;
                       end 
                      
                  10'sd362/*362:xpc10*/:  begin 
                       xpc10 <= 10'sd355/*355:xpc10*/;
                       Tspr27_2_V_3 <= (-64'sh20_0000_0000_0000<$signed((Tspr27_2_V_1<<32'sd1)));
                       end 
                      
                  10'sd363/*363:xpc10*/:  begin 
                       xpc10 <= 10'sd245/*245:xpc10*/;
                       Tdsi3_5_V_2 <= 32'sd1+Tdsi3_5_V_2;
                       Tdsi3_5_V_0 <= Tsf1SPILL12_256;
                       end 
                      
                  10'sd365/*365:xpc10*/:  begin 
                       xpc10 <= 10'sd366/*366:xpc10*/;
                       Tssu2_4_V_4 <= 64'sh_4000_0000_0000_0000|Tssu2_4_V_4;
                       end 
                      
                  10'sd366/*366:xpc10*/:  begin 
                       xpc10 <= 10'sd367/*367:xpc10*/;
                       Tssu2_4_V_6 <= Tssu2_4_V_4+(0-Tssu2_4_V_5);
                       end 
                      
                  10'sd367/*367:xpc10*/:  begin 
                       xpc10 <= 10'sd368/*368:xpc10*/;
                       Tssu2_4_V_3 <= rtl_signed_bitextract0(-16'sd1+rtl_signed_bitextract0(Tssu2_4_V_1));
                       end 
                      
                  10'sd368/*368:xpc10*/:  begin 
                       xpc10 <= 10'sd369/*369:xpc10*/;
                       Tsco0_2_V_1 <= 8'h0;
                       Tsco0_2_V_0 <= Tssu2_4_V_6;
                       end 
                      
                  10'sd372/*372:xpc10*/:  begin 
                       xpc10 <= 10'sd373/*373:xpc10*/;
                       Tsco3_7_V_0 <= (Tsco3_7_V_0<<32'sd8);
                       end 
                      
                  10'sd373/*373:xpc10*/:  begin 
                       xpc10 <= 10'sd374/*374:xpc10*/;
                       Tsco3_7_V_1 <= rtl_unsigned_bitextract3(Tsco3_7_V_1+A_8_US_CC_SCALbx14_ARA0[$unsigned((Tsco3_7_V_0>>32'sd24))]
                      );

                       end 
                      
                  10'sd374/*374:xpc10*/:  begin 
                       xpc10 <= 10'sd375/*375:xpc10*/;
                       Tsco0_2_V_1 <= rtl_unsigned_bitextract3(Tsco0_2_V_1+Tsco3_7_V_1);
                       end 
                      
                  10'sd375/*375:xpc10*/:  begin 
                       xpc10 <= 10'sd376/*376:xpc10*/;
                       Tsno34_9_V_0 <= $unsigned(-32'sd1+rtl_sign_extend10(Tsco0_2_V_1));
                       end 
                      
                  10'sd376/*376:xpc10*/:  begin 
                       xpc10 <= 10'sd377/*377:xpc10*/;
                       Tsro0_16_V_0 <= rtl_signed_bitextract0(rtl_sign_extend2(Tssu2_4_V_3)+(0-Tsno34_9_V_0));
                       end 
                      
                  10'sd377/*377:xpc10*/:  begin 
                       xpc10 <= 10'sd378/*378:xpc10*/;
                       Tsro0_16_V_1 <= (Tssu2_4_V_6<<(32'sd63&Tsno34_9_V_0));
                       end 
                      
                  10'sd379/*379:xpc10*/:  begin 
                       xpc10 <= 10'sd380/*380:xpc10*/;
                       Tsro0_16_V_6 <= rtl_signed_bitextract9(64'sh3ff&Tsro0_16_V_1);
                       Tsro0_16_V_5 <= 16'sh200;
                       end 
                      
                  10'sd382/*382:xpc10*/:  begin 
                       xpc10 <= 10'sd383/*383:xpc10*/;
                       Tsr0_SPILL_256 <= fastspilldup72;
                       Tsr0_SPILL_260 <= fastspilldup72;
                       end 
                      
                  10'sd384/*384:xpc10*/:  begin 
                       xpc10 <= 10'sd385/*385:xpc10*/;
                       Tsr0_SPILL_259 <= Tsr0_SPILL_257+(0-Tsr0_SPILL_258);
                       end 
                      
                  10'sd385/*385:xpc10*/:  begin 
                       xpc10 <= 10'sd363/*363:xpc10*/;
                       Tsf1SPILL12_256 <= Tsr0_SPILL_259;
                       Tss2_SPILL_256 <= Tsr0_SPILL_259;
                       end 
                      
                  10'sd386/*386:xpc10*/:  begin 
                       xpc10 <= 10'sd385/*385:xpc10*/;
                       Tsr0_SPILL_259 <= Tsr0_SPILL_257+(0-Tsr0_SPILL_258);
                       end 
                      
                  10'sd387/*387:xpc10*/:  begin 
                       xpc10 <= 10'sd388/*388:xpc10*/;
                       Tsro0_16_V_0 <= 16'sh0;
                       Tsro0_16_V_1 <= Tssh18_7_V_0;
                       end 
                      
                  10'sd388/*388:xpc10*/:  begin 
                       xpc10 <= 10'sd389/*389:xpc10*/;
                       Tsro0_16_V_6 <= rtl_signed_bitextract9(64'sh3ff&Tsro0_16_V_1);
                       end 
                      
                  10'sd391/*391:xpc10*/:  begin 
                       xpc10 <= 10'sd392/*392:xpc10*/;
                       Tsro0_16_V_1 <= (Tsro0_16_V_1+rtl_sign_extend4(Tsro0_16_V_5)>>32'sd10);
                       end 
                      
                  10'sd394/*394:xpc10*/:  begin 
                       xpc10 <= 10'sd395/*395:xpc10*/;
                       Tsr0_SPILL_259 <= Tsro0_16_V_1+(Tsp27_SPILL_256<<32'sd63)+(rtl_sign_extend4(Tsro0_16_V_0)<<32'sd52);
                       end 
                      
                  10'sd395/*395:xpc10*/:  begin 
                       xpc10 <= 10'sd363/*363:xpc10*/;
                       Tsf1SPILL12_256 <= Tsr0_SPILL_259;
                       Tss2_SPILL_256 <= Tsr0_SPILL_259;
                       end 
                      
                  10'sd396/*396:xpc10*/:  begin 
                       xpc10 <= 10'sd395/*395:xpc10*/;
                       Tsr0_SPILL_259 <= Tsro0_16_V_1+(Tsp27_SPILL_256<<32'sd63)+(rtl_sign_extend4(Tsro0_16_V_0)<<32'sd52);
                       end 
                      
                  10'sd397/*397:xpc10*/:  begin 
                       xpc10 <= 10'sd398/*398:xpc10*/;
                       Tss18_SPILL_256 <= fastspilldup74;
                       Tss18_SPILL_259 <= fastspilldup74;
                       end 
                      
                  10'sd399/*399:xpc10*/:  begin 
                       xpc10 <= 10'sd400/*400:xpc10*/;
                       Tssh18_7_V_0 <= Tss18_SPILL_258|Tss18_SPILL_257;
                       end 
                      
                  10'sd400/*400:xpc10*/:  begin 
                       xpc10 <= 10'sd388/*388:xpc10*/;
                       Tsro0_16_V_0 <= 16'sh0;
                       Tsro0_16_V_1 <= Tssh18_7_V_0;
                       end 
                      
                  10'sd401/*401:xpc10*/:  begin 
                       xpc10 <= 10'sd400/*400:xpc10*/;
                       Tssh18_7_V_0 <= Tss18_SPILL_258|Tss18_SPILL_257;
                       end 
                      
                  10'sd402/*402:xpc10*/:  begin 
                       xpc10 <= 10'sd403/*403:xpc10*/;
                       Tsro0_16_V_1 <= Tss18_SPILL_260;
                       Tssh18_7_V_0 <= Tss18_SPILL_260;
                       end 
                      
                  10'sd403/*403:xpc10*/:  begin 
                       xpc10 <= 10'sd389/*389:xpc10*/;
                       Tsro0_16_V_6 <= rtl_signed_bitextract9(64'sh3ff&Tsro0_16_V_1);
                       Tsro0_16_V_0 <= 16'sh0;
                       end 
                      
                  10'sd404/*404:xpc10*/:  begin 
                       xpc10 <= 10'sd403/*403:xpc10*/;
                       Tsro0_16_V_1 <= Tss18_SPILL_260;
                       Tssh18_7_V_0 <= Tss18_SPILL_260;
                       end 
                      
                  10'sd405/*405:xpc10*/:  begin 
                       xpc10 <= 10'sd370/*370:xpc10*/;
                       Tsco3_7_V_0 <= rtl_unsigned_bitextract1(64'h_ffff_ffff&Tsco0_2_V_0);
                       end 
                      
                  10'sd406/*406:xpc10*/:  begin 
                       xpc10 <= 10'sd407/*407:xpc10*/;
                       Tss32_SPILL_256 <= fastspilldup70;
                       Tss32_SPILL_259 <= fastspilldup70;
                       end 
                      
                  10'sd408/*408:xpc10*/:  begin 
                       xpc10 <= 10'sd409/*409:xpc10*/;
                       Tssh32_5_V_0 <= Tss32_SPILL_258|Tss32_SPILL_257;
                       end 
                      
                  10'sd409/*409:xpc10*/:  begin 
                       xpc10 <= 10'sd366/*366:xpc10*/;
                       Tssu2_4_V_4 <= 64'sh_4000_0000_0000_0000|Tssu2_4_V_4;
                       Tssu2_4_V_5 <= Tssh32_5_V_0;
                       end 
                      
                  10'sd410/*410:xpc10*/:  begin 
                       xpc10 <= 10'sd409/*409:xpc10*/;
                       Tssh32_5_V_0 <= Tss32_SPILL_258|Tss32_SPILL_257;
                       end 
                      
                  10'sd411/*411:xpc10*/:  begin 
                       xpc10 <= 10'sd366/*366:xpc10*/;
                       Tssu2_4_V_4 <= 64'sh_4000_0000_0000_0000|Tssu2_4_V_4;
                       Tssu2_4_V_5 <= Tssh32_5_V_0;
                       end 
                      
                  10'sd414/*414:xpc10*/:  begin 
                       xpc10 <= 10'sd415/*415:xpc10*/;
                       Tspr18_2_V_3 <= (-64'sh20_0000_0000_0000<$signed((Tspr18_2_V_1<<32'sd1)));
                       Tspr18_2_V_2 <= rtl_unsigned_bitextract5(Tsf0SPILL10_256);
                       end 
                      
                  10'sd416/*416:xpc10*/:  begin 
                       xpc10 <= 10'sd417/*417:xpc10*/;
                       Tspr18_2_V_0 <= 64'sh8_0000_0000_0000|Tspr18_2_V_0;
                       Tspr18_2_V_4 <= rtl_unsigned_bitextract5(Tsf0SPILL12_256);
                       end 
                      
                  10'sd417/*417:xpc10*/:  begin 
                       xpc10 <= 10'sd418/*418:xpc10*/;
                       Tspr18_2_V_1 <= 64'sh8_0000_0000_0000|Tspr18_2_V_1;
                       end 
                      
                  10'sd420/*420:xpc10*/:  begin 
                       xpc10 <= 10'sd244/*244:xpc10*/;
                       Tdsi3_5_V_0 <= Tss2_SPILL_256;
                       Tsf1SPILL12_256 <= Tss2_SPILL_256;
                       end 
                      
                  10'sd421/*421:xpc10*/:  begin 
                       xpc10 <= 10'sd417/*417:xpc10*/;
                       Tspr18_2_V_0 <= 64'sh8_0000_0000_0000|Tspr18_2_V_0;
                       end 
                      
                  10'sd422/*422:xpc10*/:  begin 
                       xpc10 <= 10'sd415/*415:xpc10*/;
                       Tspr18_2_V_3 <= (-64'sh20_0000_0000_0000<$signed((Tspr18_2_V_1<<32'sd1)));
                       end 
                      
                  10'sd423/*423:xpc10*/:  begin 
                       xpc10 <= 10'sd244/*244:xpc10*/;
                       Tdsi3_5_V_0 <= Tss2_SPILL_256;
                       Tsf1SPILL12_256 <= Tss2_SPILL_256;
                       end 
                      
                  10'sd425/*425:xpc10*/:  begin 
                       xpc10 <= 10'sd426/*426:xpc10*/;
                       Tssu2_4_V_5 <= 64'sh_4000_0000_0000_0000|Tssu2_4_V_5;
                       end 
                      
                  10'sd426/*426:xpc10*/:  begin 
                       xpc10 <= 10'sd427/*427:xpc10*/;
                       Tssu2_4_V_6 <= Tssu2_4_V_5+(0-Tssu2_4_V_4);
                       end 
                      
                  10'sd427/*427:xpc10*/:  begin 
                       xpc10 <= 10'sd428/*428:xpc10*/;
                       Tssu2_4_V_0 <= (Tssu2_4_V_0==32'sd0/*0:Tssu2.4_V_0*/);
                       Tssu2_4_V_3 <= rtl_signed_bitextract0(Tssu2_4_V_2);
                       end 
                      
                  10'sd428/*428:xpc10*/:  begin 
                       xpc10 <= 10'sd368/*368:xpc10*/;
                       Tssu2_4_V_3 <= rtl_signed_bitextract0(-16'sd1+Tssu2_4_V_3);
                       end 
                      
                  10'sd429/*429:xpc10*/:  begin 
                       xpc10 <= 10'sd430/*430:xpc10*/;
                       Tss23_SPILL_256 <= fastspilldup68;
                       Tss23_SPILL_259 <= fastspilldup68;
                       end 
                      
                  10'sd431/*431:xpc10*/:  begin 
                       xpc10 <= 10'sd432/*432:xpc10*/;
                       Tssh23_6_V_0 <= Tss23_SPILL_258|Tss23_SPILL_257;
                       end 
                      
                  10'sd432/*432:xpc10*/:  begin 
                       xpc10 <= 10'sd426/*426:xpc10*/;
                       Tssu2_4_V_5 <= 64'sh_4000_0000_0000_0000|Tssu2_4_V_5;
                       Tssu2_4_V_4 <= Tssh23_6_V_0;
                       end 
                      
                  10'sd433/*433:xpc10*/:  begin 
                       xpc10 <= 10'sd432/*432:xpc10*/;
                       Tssh23_6_V_0 <= Tss23_SPILL_258|Tss23_SPILL_257;
                       end 
                      
                  10'sd434/*434:xpc10*/:  begin 
                       xpc10 <= 10'sd426/*426:xpc10*/;
                       Tssu2_4_V_5 <= 64'sh_4000_0000_0000_0000|Tssu2_4_V_5;
                       Tssu2_4_V_4 <= Tssh23_6_V_0;
                       end 
                      
                  10'sd437/*437:xpc10*/:  begin 
                       xpc10 <= 10'sd438/*438:xpc10*/;
                       Tspr7_3_V_3 <= (-64'sh20_0000_0000_0000<$signed((Tspr7_3_V_1<<32'sd1)));
                       Tspr7_3_V_2 <= rtl_unsigned_bitextract5(Tsf0SPILL10_256);
                       end 
                      
                  10'sd439/*439:xpc10*/:  begin 
                       xpc10 <= 10'sd440/*440:xpc10*/;
                       Tspr7_3_V_0 <= 64'sh8_0000_0000_0000|Tspr7_3_V_0;
                       Tspr7_3_V_4 <= rtl_unsigned_bitextract5(Tsf0SPILL12_256);
                       end 
                      
                  10'sd440/*440:xpc10*/:  begin 
                       xpc10 <= 10'sd441/*441:xpc10*/;
                       Tspr7_3_V_1 <= 64'sh8_0000_0000_0000|Tspr7_3_V_1;
                       end 
                      
                  10'sd443/*443:xpc10*/:  begin 
                       xpc10 <= 10'sd244/*244:xpc10*/;
                       Tdsi3_5_V_0 <= Tss2_SPILL_256;
                       Tsf1SPILL12_256 <= Tss2_SPILL_256;
                       end 
                      
                  10'sd444/*444:xpc10*/:  begin 
                       xpc10 <= 10'sd440/*440:xpc10*/;
                       Tspr7_3_V_0 <= 64'sh8_0000_0000_0000|Tspr7_3_V_0;
                       end 
                      
                  10'sd445/*445:xpc10*/:  begin 
                       xpc10 <= 10'sd438/*438:xpc10*/;
                       Tspr7_3_V_3 <= (-64'sh20_0000_0000_0000<$signed((Tspr7_3_V_1<<32'sd1)));
                       end 
                      
                  10'sd446/*446:xpc10*/:  begin 
                       xpc10 <= 10'sd363/*363:xpc10*/;
                       Tsf1SPILL12_256 <= 64'h_7fff_ffff_ffff_ffff;
                       Tss2_SPILL_256 <= 64'h_7fff_ffff_ffff_ffff;
                       end 
                      
                  10'sd448/*448:xpc10*/:  begin 
                       xpc10 <= 10'sd244/*244:xpc10*/;
                       Tdsi3_5_V_0 <= Tss2_SPILL_256;
                       Tsf1SPILL12_256 <= Tss2_SPILL_256;
                       end 
                      
                  10'sd451/*451:xpc10*/:  begin 
                       xpc10 <= 10'sd223/*223:xpc10*/;
                       Tspr2_2_V_0 <= 64'sh8_0000_0000_0000|Tspr2_2_V_0;
                       end 
                      
                  10'sd452/*452:xpc10*/:  begin 
                       xpc10 <= 10'sd221/*221:xpc10*/;
                       Tspr2_2_V_3 <= (-64'sh20_0000_0000_0000<$signed((Tspr2_2_V_1<<32'sd1)));
                       end 
                      
                  10'sd454/*454:xpc10*/:  begin 
                       xpc10 <= 10'sd455/*455:xpc10*/;
                       Tspr5_2_V_3 <= (-64'sh20_0000_0000_0000<$signed((Tspr5_2_V_1<<32'sd1)));
                       Tspr5_2_V_2 <= rtl_unsigned_bitextract5(Tsf0SPILL10_256);
                       end 
                      
                  10'sd456/*456:xpc10*/:  begin 
                       xpc10 <= 10'sd457/*457:xpc10*/;
                       Tspr5_2_V_0 <= 64'sh8_0000_0000_0000|Tspr5_2_V_0;
                       Tspr5_2_V_4 <= rtl_unsigned_bitextract5(Tsf0SPILL12_256);
                       end 
                      
                  10'sd457/*457:xpc10*/:  begin 
                       xpc10 <= 10'sd458/*458:xpc10*/;
                       Tspr5_2_V_1 <= 64'sh8_0000_0000_0000|Tspr5_2_V_1;
                       end 
                      
                  10'sd461/*461:xpc10*/:  begin 
                       xpc10 <= 10'sd457/*457:xpc10*/;
                       Tspr5_2_V_0 <= 64'sh8_0000_0000_0000|Tspr5_2_V_0;
                       end 
                      
                  10'sd462/*462:xpc10*/:  begin 
                       xpc10 <= 10'sd455/*455:xpc10*/;
                       Tspr5_2_V_3 <= (-64'sh20_0000_0000_0000<$signed((Tspr5_2_V_1<<32'sd1)));
                       end 
                      
                  10'sd463/*463:xpc10*/:  begin 
                       xpc10 <= 10'sd464/*464:xpc10*/;
                       Tdsi3_5_V_1 <= 64'h_7fff_ffff_ffff_ffff;
                       Tsf1SPILL10_256 <= 64'h_7fff_ffff_ffff_ffff;
                       end 
                      
                  10'sd469/*469:xpc10*/:  begin 
                       xpc10 <= 10'sd470/*470:xpc10*/;
                       Tspr10_2_V_3 <= (-64'sh20_0000_0000_0000<$signed((Tspr10_2_V_1<<32'sd1)));
                       Tspr10_2_V_2 <= rtl_unsigned_bitextract5(Tsf0SPILL10_256);
                       end 
                      
                  10'sd471/*471:xpc10*/:  begin 
                       xpc10 <= 10'sd472/*472:xpc10*/;
                       Tspr10_2_V_0 <= 64'sh8_0000_0000_0000|Tspr10_2_V_0;
                       Tspr10_2_V_4 <= rtl_unsigned_bitextract5(Tsf0SPILL12_256);
                       end 
                      
                  10'sd472/*472:xpc10*/:  begin 
                       xpc10 <= 10'sd473/*473:xpc10*/;
                       Tspr10_2_V_1 <= 64'sh8_0000_0000_0000|Tspr10_2_V_1;
                       end 
                      
                  10'sd476/*476:xpc10*/:  begin 
                       xpc10 <= 10'sd472/*472:xpc10*/;
                       Tspr10_2_V_0 <= 64'sh8_0000_0000_0000|Tspr10_2_V_0;
                       end 
                      
                  10'sd477/*477:xpc10*/:  begin 
                       xpc10 <= 10'sd470/*470:xpc10*/;
                       Tspr10_2_V_3 <= (-64'sh20_0000_0000_0000<$signed((Tspr10_2_V_1<<32'sd1)));
                       end 
                      
                  10'sd479/*479:xpc10*/:  begin 
                       xpc10 <= 10'sd464/*464:xpc10*/;
                       Tdsi3_5_V_1 <= 64'h_7fff_ffff_ffff_ffff;
                       Tsf1SPILL10_256 <= 64'h_7fff_ffff_ffff_ffff;
                       end 
                      
                  10'sd485/*485:xpc10*/:  begin 
                       xpc10 <= 10'sd486/*486:xpc10*/;
                       Tsco3_7_V_0 <= (Tsco3_7_V_0<<32'sd8);
                       end 
                      
                  10'sd486/*486:xpc10*/:  begin 
                       xpc10 <= 10'sd487/*487:xpc10*/;
                       Tsco3_7_V_1 <= rtl_unsigned_bitextract3(Tsco3_7_V_1+A_8_US_CC_SCALbx14_ARA0[$unsigned((Tsco3_7_V_0>>32'sd24))]
                      );

                       end 
                      
                  10'sd487/*487:xpc10*/:  begin 
                       xpc10 <= 10'sd488/*488:xpc10*/;
                       Tsco0_2_V_1 <= rtl_unsigned_bitextract3(Tsco0_2_V_1+Tsco3_7_V_1);
                       end 
                      
                  10'sd488/*488:xpc10*/:  begin 
                       xpc10 <= 10'sd489/*489:xpc10*/;
                       Tsno18_4_V_0 <= $unsigned(-32'sd11+rtl_sign_extend10(Tsco0_2_V_1));
                       end 
                      
                  10'sd489/*489:xpc10*/:  begin 
                       xpc10 <= 10'sd490/*490:xpc10*/;
                       Tsfl1_18_V_7 <= (Tsfl1_18_V_7<<(32'sd63&Tsno18_4_V_0));
                       end 
                      
                  10'sd490/*490:xpc10*/:  begin 
                       xpc10 <= 10'sd491/*491:xpc10*/;
                       Tsfl1_18_V_4 <= rtl_signed_bitextract0(rtl_sign_extend2(16'sd1)+(0-Tsno18_4_V_0));
                       end 
                      
                  10'sd496/*496:xpc10*/:  begin 
                       xpc10 <= 10'sd497/*497:xpc10*/;
                       Tsco3_7_V_0 <= (Tsco3_7_V_0<<32'sd8);
                       end 
                      
                  10'sd497/*497:xpc10*/:  begin 
                       xpc10 <= 10'sd498/*498:xpc10*/;
                       Tsco3_7_V_1 <= rtl_unsigned_bitextract3(Tsco3_7_V_1+A_8_US_CC_SCALbx14_ARA0[$unsigned((Tsco3_7_V_0>>32'sd24))]
                      );

                       end 
                      
                  10'sd498/*498:xpc10*/:  begin 
                       xpc10 <= 10'sd499/*499:xpc10*/;
                       Tsco0_2_V_1 <= rtl_unsigned_bitextract3(Tsco0_2_V_1+Tsco3_7_V_1);
                       end 
                      
                  10'sd499/*499:xpc10*/:  begin 
                       xpc10 <= 10'sd500/*500:xpc10*/;
                       Tsno22_4_V_0 <= $unsigned(-32'sd11+rtl_sign_extend10(Tsco0_2_V_1));
                       end 
                      
                  10'sd500/*500:xpc10*/:  begin 
                       xpc10 <= 10'sd501/*501:xpc10*/;
                       Tsfl1_18_V_6 <= (Tsfl1_18_V_6<<(32'sd63&Tsno22_4_V_0));
                       end 
                      
                  10'sd501/*501:xpc10*/:  begin 
                       xpc10 <= 10'sd502/*502:xpc10*/;
                       Tsfl1_18_V_3 <= rtl_signed_bitextract0(rtl_sign_extend2(16'sd1)+(0-Tsno22_4_V_0));
                       end 
                      
                  10'sd502/*502:xpc10*/:  begin 
                       xpc10 <= 10'sd503/*503:xpc10*/;
                       Tsfl1_18_V_5 <= rtl_signed_bitextract0(rtl_sign_extend2(16'sd1021)+rtl_sign_extend2(Tsfl1_18_V_3)+(0-Tsfl1_18_V_4
                      ));

                       end 
                      
                  10'sd503/*503:xpc10*/:  begin 
                       xpc10 <= 10'sd504/*504:xpc10*/;
                       Tsfl1_18_V_6 <= ((64'sh10_0000_0000_0000|Tsfl1_18_V_6)<<32'sd10);
                       end 
                      
                  10'sd504/*504:xpc10*/:  begin 
                       xpc10 <= 10'sd505/*505:xpc10*/;
                       Tsfl1_18_V_7 <= ((64'sh10_0000_0000_0000|Tsfl1_18_V_7)<<32'sd11);
                       end 
                      
                  10'sd506/*506:xpc10*/:  begin 
                       xpc10 <= 10'sd507/*507:xpc10*/;
                       Tsfl1_18_V_5 <= rtl_signed_bitextract0(16'sd1+Tsfl1_18_V_5);
                       end 
                      
                  10'sd509/*509:xpc10*/:  begin 
                       xpc10 <= 10'sd510/*510:xpc10*/;
                       Tsmu26_4_V_0 <= rtl_unsigned_bitextract1((Tsfl1_18_V_7>>32'sd32));
                       end 
                      
                  10'sd510/*510:xpc10*/:  begin 
                       xpc10 <= 10'sd511/*511:xpc10*/;
                       Tsmu26_4_V_3 <= rtl_unsigned_bitextract1(64'h_ffff_ffff&Tsfl1_18_V_8);
                       end 
                      
                  10'sd511/*511:xpc10*/:  begin 
                       xpc10 <= 10'sd512/*512:xpc10*/;
                       Tsmu26_4_V_2 <= rtl_unsigned_bitextract1((Tsfl1_18_V_8>>32'sd32));
                       end 
                      
                  10'sd512/*512:xpc10*/:  begin 
                       xpc10 <= 10'sd513/*513:xpc10*/;
                       Tsmu26_4_V_7 <= rtl_unsigned_extend7(Tsmu26_4_V_1)*rtl_unsigned_extend7(Tsmu26_4_V_3);
                       end 
                      
                  10'sd513/*513:xpc10*/:  begin 
                       xpc10 <= 10'sd514/*514:xpc10*/;
                       Tsmu26_4_V_5 <= rtl_unsigned_extend7(Tsmu26_4_V_1)*rtl_unsigned_extend7(Tsmu26_4_V_2);
                       end 
                      
                  10'sd514/*514:xpc10*/:  begin 
                       xpc10 <= 10'sd515/*515:xpc10*/;
                       Tsmu26_4_V_6 <= rtl_unsigned_extend7(Tsmu26_4_V_0)*rtl_unsigned_extend7(Tsmu26_4_V_3);
                       end 
                      
                  10'sd515/*515:xpc10*/:  begin 
                       xpc10 <= 10'sd516/*516:xpc10*/;
                       Tsmu26_4_V_4 <= rtl_unsigned_extend7(Tsmu26_4_V_0)*rtl_unsigned_extend7(Tsmu26_4_V_2);
                       end 
                      
                  10'sd516/*516:xpc10*/:  begin 
                       xpc10 <= 10'sd517/*517:xpc10*/;
                       Tsmu26_4_V_5 <= Tsmu26_4_V_5+Tsmu26_4_V_6;
                       end 
                      
                  10'sd518/*518:xpc10*/:  begin 
                       xpc10 <= 10'sd519/*519:xpc10*/;
                       Tsm26_SPILL_264 <= Tsmu26_4_V_4;
                       fastspilldup46 <= Tsmu26_4_V_4;
                       end 
                      
                  10'sd520/*520:xpc10*/:  begin 
                       xpc10 <= 10'sd521/*521:xpc10*/;
                       Tsmu26_4_V_4 <= Tsm26_SPILL_257+(Tsm26_SPILL_259<<32'sd32)+(Tsmu26_4_V_5>>32'sd32);
                       end 
                      
                  10'sd521/*521:xpc10*/:  begin 
                       xpc10 <= 10'sd522/*522:xpc10*/;
                       Tsmu26_4_V_5 <= (Tsmu26_4_V_5<<32'sd32);
                       end 
                      
                  10'sd522/*522:xpc10*/:  begin 
                       xpc10 <= 10'sd523/*523:xpc10*/;
                       Tsmu26_4_V_7 <= Tsmu26_4_V_7+Tsmu26_4_V_5;
                       end 
                      
                  10'sd523/*523:xpc10*/:  begin 
                       xpc10 <= 10'sd524/*524:xpc10*/;
                       Tsm26_SPILL_263 <= Tsmu26_4_V_4;
                       fastspilldup48 <= Tsmu26_4_V_4;
                       end 
                      
                  10'sd525/*525:xpc10*/:  begin 
                       xpc10 <= 10'sd526/*526:xpc10*/;
                       Tsmu26_4_V_4 <= Tsm26_SPILL_260+Tsm26_SPILL_262;
                       end 
                      
                  10'sd526/*526:xpc10*/:  begin 
                       xpc10 <= 10'sd527/*527:xpc10*/;
                       Tsfl1_18_V_11 <= Tsmu26_4_V_4;
                       Tsfl1_18_V_12 <= Tsmu26_4_V_7;
                       end 
                      
                  10'sd527/*527:xpc10*/:  begin 
                       xpc10 <= 10'sd528/*528:xpc10*/;
                       Tsfl1_18_V_10 <= 64'sh0+(0-Tsfl1_18_V_12);
                       end 
                      
                  10'sd528/*528:xpc10*/:  begin 
                       xpc10 <= 10'sd529/*529:xpc10*/;
                       fastspilldup50 <= Tsfl1_18_V_6+(0-Tsfl1_18_V_11);
                       end 
                      
                  10'sd529/*529:xpc10*/:  begin 
                       xpc10 <= 10'sd530/*530:xpc10*/;
                       Tss26_SPILL_257 <= fastspilldup50;
                       Tss26_SPILL_262 <= fastspilldup50;
                       end 
                      
                  10'sd531/*531:xpc10*/:  begin 
                       xpc10 <= 10'sd532/*532:xpc10*/;
                       Tsfl1_18_V_9 <= Tss26_SPILL_259+(0-Tss26_SPILL_260);
                       end 
                      
                  10'sd534/*534:xpc10*/:  begin 
                       xpc10 <= 10'sd535/*535:xpc10*/;
                       Tsfl1_18_V_8 <= Tsf1SPILL10_257|Tsf1SPILL10_259;
                       end 
                      
                  10'sd535/*535:xpc10*/:  begin 
                       xpc10 <= 10'sd536/*536:xpc10*/;
                       Tsro33_4_V_1 <= Tsfl1_18_V_8;
                       Tsro33_4_V_0 <= rtl_signed_bitextract0(Tsfl1_18_V_5);
                       end 
                      
                  10'sd537/*537:xpc10*/:  begin 
                       xpc10 <= 10'sd538/*538:xpc10*/;
                       Tsro33_4_V_6 <= rtl_signed_bitextract9(64'sh3ff&Tsro33_4_V_1);
                       Tsro33_4_V_5 <= 16'sh200;
                       end 
                      
                  10'sd540/*540:xpc10*/:  begin 
                       xpc10 <= 10'sd541/*541:xpc10*/;
                       Tsr33_SPILL_256 <= fastspilldup56;
                       Tsr33_SPILL_260 <= fastspilldup56;
                       end 
                      
                  10'sd542/*542:xpc10*/:  begin 
                       xpc10 <= 10'sd543/*543:xpc10*/;
                       Tsr33_SPILL_259 <= Tsr33_SPILL_257+(0-Tsr33_SPILL_258);
                       end 
                      
                  10'sd543/*543:xpc10*/:  begin 
                       xpc10 <= 10'sd464/*464:xpc10*/;
                       Tdsi3_5_V_1 <= Tsr33_SPILL_259;
                       Tsf1SPILL10_256 <= Tsr33_SPILL_259;
                       end 
                      
                  10'sd544/*544:xpc10*/:  begin 
                       xpc10 <= 10'sd543/*543:xpc10*/;
                       Tsr33_SPILL_259 <= Tsr33_SPILL_257+(0-Tsr33_SPILL_258);
                       end 
                      
                  10'sd545/*545:xpc10*/:  begin 
                       xpc10 <= 10'sd546/*546:xpc10*/;
                       Tsro33_4_V_0 <= 16'sh0;
                       Tsro33_4_V_1 <= Tssh18_7_V_0;
                       end 
                      
                  10'sd546/*546:xpc10*/:  begin 
                       xpc10 <= 10'sd547/*547:xpc10*/;
                       Tsro33_4_V_6 <= rtl_signed_bitextract9(64'sh3ff&Tsro33_4_V_1);
                       end 
                      
                  10'sd549/*549:xpc10*/:  begin 
                       xpc10 <= 10'sd550/*550:xpc10*/;
                       Tsro33_4_V_1 <= (Tsro33_4_V_1+rtl_sign_extend4(Tsro33_4_V_5)>>32'sd10);
                       end 
                      
                  10'sd552/*552:xpc10*/:  begin 
                       xpc10 <= 10'sd553/*553:xpc10*/;
                       Tsr33_SPILL_259 <= Tsro33_4_V_1+(Tsp27_SPILL_256<<32'sd63)+(rtl_sign_extend4(Tsro33_4_V_0)<<32'sd52);
                       end 
                      
                  10'sd553/*553:xpc10*/:  begin 
                       xpc10 <= 10'sd464/*464:xpc10*/;
                       Tdsi3_5_V_1 <= Tsr33_SPILL_259;
                       Tsf1SPILL10_256 <= Tsr33_SPILL_259;
                       end 
                      
                  10'sd554/*554:xpc10*/:  begin 
                       xpc10 <= 10'sd553/*553:xpc10*/;
                       Tsr33_SPILL_259 <= Tsro33_4_V_1+(Tsp27_SPILL_256<<32'sd63)+(rtl_sign_extend4(Tsro33_4_V_0)<<32'sd52);
                       end 
                      
                  10'sd555/*555:xpc10*/:  begin 
                       xpc10 <= 10'sd556/*556:xpc10*/;
                       Tss18_SPILL_256 <= fastspilldup58;
                       Tss18_SPILL_259 <= fastspilldup58;
                       end 
                      
                  10'sd557/*557:xpc10*/:  begin 
                       xpc10 <= 10'sd558/*558:xpc10*/;
                       Tssh18_7_V_0 <= Tss18_SPILL_258|Tss18_SPILL_257;
                       end 
                      
                  10'sd558/*558:xpc10*/:  begin 
                       xpc10 <= 10'sd546/*546:xpc10*/;
                       Tsro33_4_V_0 <= 16'sh0;
                       Tsro33_4_V_1 <= Tssh18_7_V_0;
                       end 
                      
                  10'sd559/*559:xpc10*/:  begin 
                       xpc10 <= 10'sd558/*558:xpc10*/;
                       Tssh18_7_V_0 <= Tss18_SPILL_258|Tss18_SPILL_257;
                       end 
                      
                  10'sd560/*560:xpc10*/:  begin 
                       xpc10 <= 10'sd561/*561:xpc10*/;
                       Tsro33_4_V_1 <= Tss18_SPILL_260;
                       Tssh18_7_V_0 <= Tss18_SPILL_260;
                       end 
                      
                  10'sd561/*561:xpc10*/:  begin 
                       xpc10 <= 10'sd547/*547:xpc10*/;
                       Tsro33_4_V_6 <= rtl_signed_bitextract9(64'sh3ff&Tsro33_4_V_1);
                       Tsro33_4_V_0 <= 16'sh0;
                       end 
                      
                  10'sd562/*562:xpc10*/:  begin 
                       xpc10 <= 10'sd561/*561:xpc10*/;
                       Tsro33_4_V_1 <= Tss18_SPILL_260;
                       Tssh18_7_V_0 <= Tss18_SPILL_260;
                       end 
                      
                  10'sd563/*563:xpc10*/:  begin 
                       xpc10 <= 10'sd535/*535:xpc10*/;
                       Tsfl1_18_V_8 <= Tsf1SPILL10_260|Tsf1SPILL10_259;
                       end 
                      
                  10'sd564/*564:xpc10*/:  begin 
                       xpc10 <= 10'sd565/*565:xpc10*/;
                       Tsad27_13_V_0 <= Tsfl1_18_V_7+Tsfl1_18_V_10;
                       end 
                      
                  10'sd565/*565:xpc10*/:  begin 
                       xpc10 <= 10'sd566/*566:xpc10*/;
                       fastspilldup52 <= 64'sh0+Tsfl1_18_V_9;
                       Tsfl1_18_V_10 <= Tsad27_13_V_0;
                       end 
                      
                  10'sd566/*566:xpc10*/:  begin 
                       xpc10 <= 10'sd567/*567:xpc10*/;
                       Tsa27_SPILL_257 <= fastspilldup52;
                       Tsa27_SPILL_262 <= fastspilldup52;
                       end 
                      
                  10'sd568/*568:xpc10*/:  begin 
                       xpc10 <= 10'sd569/*569:xpc10*/;
                       Tsfl1_18_V_9 <= Tsa27_SPILL_260+Tsa27_SPILL_259;
                       end 
                      
                  10'sd570/*570:xpc10*/:  begin 
                       xpc10 <= 10'sd569/*569:xpc10*/;
                       Tsfl1_18_V_9 <= Tsa27_SPILL_260+Tsa27_SPILL_259;
                       end 
                      
                  10'sd571/*571:xpc10*/:  begin 
                       xpc10 <= 10'sd532/*532:xpc10*/;
                       Tsfl1_18_V_9 <= Tss26_SPILL_259+(0-Tss26_SPILL_260);
                       end 
                      
                  10'sd572/*572:xpc10*/:  begin 
                       xpc10 <= 10'sd526/*526:xpc10*/;
                       Tsmu26_4_V_4 <= Tsm26_SPILL_263+Tsm26_SPILL_262;
                       end 
                      
                  10'sd573/*573:xpc10*/:  begin 
                       xpc10 <= 10'sd521/*521:xpc10*/;
                       Tsmu26_4_V_4 <= Tsm26_SPILL_264+(Tsm26_SPILL_259<<32'sd32)+(Tsmu26_4_V_5>>32'sd32);
                       end 
                      
                  10'sd575/*575:xpc10*/:  begin 
                       xpc10 <= 10'sd576/*576:xpc10*/;
                       Tsmu5_7_V_1 <= rtl_unsigned_bitextract1(64'h_ffff_ffff&Tsfl1_18_V_7);
                       end 
                      
                  10'sd576/*576:xpc10*/:  begin 
                       xpc10 <= 10'sd577/*577:xpc10*/;
                       Tsmu5_7_V_0 <= rtl_unsigned_bitextract1((Tsfl1_18_V_7>>32'sd32));
                       end 
                      
                  10'sd577/*577:xpc10*/:  begin 
                       xpc10 <= 10'sd578/*578:xpc10*/;
                       Tsmu5_7_V_3 <= rtl_unsigned_bitextract1(64'h_ffff_ffff&Tses25_5_V_6);
                       end 
                      
                  10'sd578/*578:xpc10*/:  begin 
                       xpc10 <= 10'sd579/*579:xpc10*/;
                       Tsmu5_7_V_2 <= rtl_unsigned_bitextract1((Tses25_5_V_6>>32'sd32));
                       end 
                      
                  10'sd579/*579:xpc10*/:  begin 
                       xpc10 <= 10'sd580/*580:xpc10*/;
                       Tsmu5_7_V_7 <= rtl_unsigned_extend7(Tsmu5_7_V_1)*rtl_unsigned_extend7(Tsmu5_7_V_3);
                       end 
                      
                  10'sd580/*580:xpc10*/:  begin 
                       xpc10 <= 10'sd581/*581:xpc10*/;
                       Tsmu5_7_V_5 <= rtl_unsigned_extend7(Tsmu5_7_V_1)*rtl_unsigned_extend7(Tsmu5_7_V_2);
                       end 
                      
                  10'sd581/*581:xpc10*/:  begin 
                       xpc10 <= 10'sd582/*582:xpc10*/;
                       Tsmu5_7_V_6 <= rtl_unsigned_extend7(Tsmu5_7_V_0)*rtl_unsigned_extend7(Tsmu5_7_V_3);
                       end 
                      
                  10'sd582/*582:xpc10*/:  begin 
                       xpc10 <= 10'sd583/*583:xpc10*/;
                       Tsmu5_7_V_4 <= rtl_unsigned_extend7(Tsmu5_7_V_0)*rtl_unsigned_extend7(Tsmu5_7_V_2);
                       end 
                      
                  10'sd583/*583:xpc10*/:  begin 
                       xpc10 <= 10'sd584/*584:xpc10*/;
                       Tsmu5_7_V_5 <= Tsmu5_7_V_5+Tsmu5_7_V_6;
                       end 
                      
                  10'sd585/*585:xpc10*/:  begin 
                       xpc10 <= 10'sd586/*586:xpc10*/;
                       Tsm5_SPILL_264 <= Tsmu5_7_V_4;
                       fastspilldup36 <= Tsmu5_7_V_4;
                       end 
                      
                  10'sd587/*587:xpc10*/:  begin 
                       xpc10 <= 10'sd588/*588:xpc10*/;
                       Tsmu5_7_V_4 <= Tsm5_SPILL_257+(Tsm5_SPILL_259<<32'sd32)+(Tsmu5_7_V_5>>32'sd32);
                       end 
                      
                  10'sd588/*588:xpc10*/:  begin 
                       xpc10 <= 10'sd589/*589:xpc10*/;
                       Tsmu5_7_V_5 <= (Tsmu5_7_V_5<<32'sd32);
                       end 
                      
                  10'sd589/*589:xpc10*/:  begin 
                       xpc10 <= 10'sd590/*590:xpc10*/;
                       Tsmu5_7_V_7 <= Tsmu5_7_V_7+Tsmu5_7_V_5;
                       end 
                      
                  10'sd590/*590:xpc10*/:  begin 
                       xpc10 <= 10'sd591/*591:xpc10*/;
                       Tsm5_SPILL_263 <= Tsmu5_7_V_4;
                       fastspilldup38 <= Tsmu5_7_V_4;
                       end 
                      
                  10'sd592/*592:xpc10*/:  begin 
                       xpc10 <= 10'sd593/*593:xpc10*/;
                       Tsmu5_7_V_4 <= Tsm5_SPILL_260+Tsm5_SPILL_262;
                       end 
                      
                  10'sd593/*593:xpc10*/:  begin 
                       xpc10 <= 10'sd594/*594:xpc10*/;
                       Tses25_5_V_4 <= Tsmu5_7_V_4;
                       Tses25_5_V_5 <= Tsmu5_7_V_7;
                       end 
                      
                  10'sd594/*594:xpc10*/:  begin 
                       xpc10 <= 10'sd595/*595:xpc10*/;
                       Tses25_5_V_3 <= 64'sh0+(0-Tses25_5_V_5);
                       end 
                      
                  10'sd595/*595:xpc10*/:  begin 
                       xpc10 <= 10'sd596/*596:xpc10*/;
                       fastspilldup40 <= Tsfl1_18_V_6+(0-Tses25_5_V_4);
                       end 
                      
                  10'sd596/*596:xpc10*/:  begin 
                       xpc10 <= 10'sd597/*597:xpc10*/;
                       Tss5_SPILL_257 <= fastspilldup40;
                       Tss5_SPILL_262 <= fastspilldup40;
                       end 
                      
                  10'sd598/*598:xpc10*/:  begin 
                       xpc10 <= 10'sd599/*599:xpc10*/;
                       Tses25_5_V_2 <= Tss5_SPILL_259+(0-Tss5_SPILL_260);
                       end 
                      
                  10'sd600/*600:xpc10*/:  begin 
                       xpc10 <= 10'sd601/*601:xpc10*/;
                       Tse25_SPILL_261 <= Tses25_5_V_6;
                       fastspilldup44 <= Tses25_5_V_6;
                       end 
                      
                  10'sd602/*602:xpc10*/:  begin 
                       xpc10 <= 10'sd603/*603:xpc10*/;
                       Tses25_5_V_6 <= Tse25_SPILL_258|Tse25_SPILL_260;
                       end 
                      
                  10'sd603/*603:xpc10*/:  begin 
                       xpc10 <= 10'sd508/*508:xpc10*/;
                       Tsfl1_18_V_8 <= Tses25_5_V_6;
                       end 
                      
                  10'sd604/*604:xpc10*/:  begin 
                       xpc10 <= 10'sd603/*603:xpc10*/;
                       Tses25_5_V_6 <= Tse25_SPILL_261|Tse25_SPILL_260;
                       end 
                      
                  10'sd605/*605:xpc10*/:  begin 
                       xpc10 <= 10'sd606/*606:xpc10*/;
                       Tses25_5_V_1 <= (Tsfl1_18_V_7<<32'sd32);
                       end 
                      
                  10'sd606/*606:xpc10*/:  begin 
                       xpc10 <= 10'sd607/*607:xpc10*/;
                       Tsad6_15_V_0 <= Tses25_5_V_3+Tses25_5_V_1;
                       end 
                      
                  10'sd607/*607:xpc10*/:  begin 
                       xpc10 <= 10'sd608/*608:xpc10*/;
                       fastspilldup42 <= Tses25_5_V_0+Tses25_5_V_2;
                       Tses25_5_V_3 <= Tsad6_15_V_0;
                       end 
                      
                  10'sd608/*608:xpc10*/:  begin 
                       xpc10 <= 10'sd609/*609:xpc10*/;
                       Tsa6_SPILL_257 <= fastspilldup42;
                       Tsa6_SPILL_262 <= fastspilldup42;
                       end 
                      
                  10'sd610/*610:xpc10*/:  begin 
                       xpc10 <= 10'sd611/*611:xpc10*/;
                       Tses25_5_V_2 <= Tsa6_SPILL_260+Tsa6_SPILL_259;
                       end 
                      
                  10'sd612/*612:xpc10*/:  begin 
                       xpc10 <= 10'sd611/*611:xpc10*/;
                       Tses25_5_V_2 <= Tsa6_SPILL_260+Tsa6_SPILL_259;
                       end 
                      
                  10'sd613/*613:xpc10*/:  begin 
                       xpc10 <= 10'sd599/*599:xpc10*/;
                       Tses25_5_V_2 <= Tss5_SPILL_259+(0-Tss5_SPILL_260);
                       end 
                      
                  10'sd614/*614:xpc10*/:  begin 
                       xpc10 <= 10'sd593/*593:xpc10*/;
                       Tsmu5_7_V_4 <= Tsm5_SPILL_263+Tsm5_SPILL_262;
                       end 
                      
                  10'sd615/*615:xpc10*/:  begin 
                       xpc10 <= 10'sd588/*588:xpc10*/;
                       Tsmu5_7_V_4 <= Tsm5_SPILL_264+(Tsm5_SPILL_259<<32'sd32)+(Tsmu5_7_V_5>>32'sd32);
                       end 
                      
                  10'sd616/*616:xpc10*/:  begin 
                       xpc10 <= 10'sd576/*576:xpc10*/;
                       Tsmu5_7_V_1 <= rtl_unsigned_bitextract1(64'h_ffff_ffff&Tsfl1_18_V_7);
                       Tses25_5_V_6 <= Tse25_SPILL_257;
                       end 
                      
                  10'sd617/*617:xpc10*/:  begin 
                       xpc10 <= 10'sd494/*494:xpc10*/;
                       Tsco3_7_V_0 <= rtl_unsigned_bitextract1(64'h_ffff_ffff&Tsco0_2_V_0);
                       end 
                      
                  10'sd618/*618:xpc10*/:  begin 
                       xpc10 <= 10'sd483/*483:xpc10*/;
                       Tsco3_7_V_0 <= rtl_unsigned_bitextract1(64'h_ffff_ffff&Tsco0_2_V_0);
                       end 
                      
                  10'sd620/*620:xpc10*/:  begin 
                       xpc10 <= 10'sd621/*621:xpc10*/;
                       Tsco5_4_V_0 <= Tsi1_SPILL_257;
                       Tsin1_17_V_1 <= Tsi1_SPILL_257;
                       end 
                      
                  10'sd623/*623:xpc10*/:  begin 
                       xpc10 <= 10'sd624/*624:xpc10*/;
                       Tsco5_4_V_0 <= (Tsco5_4_V_0<<32'sd8);
                       end 
                      
                  10'sd624/*624:xpc10*/:  begin 
                       xpc10 <= 10'sd625/*625:xpc10*/;
                       Tsco5_4_V_1 <= rtl_unsigned_bitextract3(Tsco5_4_V_1+A_8_US_CC_SCALbx14_ARA0[$unsigned((Tsco5_4_V_0>>32'sd24))]
                      );

                       end 
                      
                  10'sd625/*625:xpc10*/:  begin 
                       xpc10 <= 10'sd626/*626:xpc10*/;
                       Tsin1_17_V_3 <= $unsigned(32'sd21+rtl_sign_extend10(Tsco5_4_V_1));
                       end 
                      
                  10'sd627/*627:xpc10*/:  begin 
                       xpc10 <= 10'sd628/*628:xpc10*/;
                       Tsi1_SPILL_256 <= (Tsp5_SPILL_256<<32'sd63)+(rtl_sign_extend11(rtl_signed_bitextract0(rtl_sign_extend2(16'sd1074
                      )+(0-Tsin1_17_V_3)))<<32'sd52)+(Tsin1_17_V_2<<(32'sd63&Tsin1_17_V_3));

                       end 
                      
                  10'sd628/*628:xpc10*/:  begin 
                       xpc10 <= 10'sd212/*212:xpc10*/;
                       Tsfl1_18_V_6 <= 64'shf_ffff_ffff_ffff&Tsf1_SPILL_256;
                       end 
                      
                  10'sd629/*629:xpc10*/:  begin 
                       xpc10 <= 10'sd628/*628:xpc10*/;
                       Tsi1_SPILL_256 <= (Tsp5_SPILL_256<<32'sd63)+(rtl_sign_extend11(rtl_signed_bitextract0(rtl_sign_extend2(16'sd1074
                      )+(0-Tsin1_17_V_3)))<<32'sd52)+(Tsin1_17_V_2<<(32'sd63&Tsin1_17_V_3));

                       end 
                      
                  10'sd630/*630:xpc10*/:  begin 
                       xpc10 <= 10'sd621/*621:xpc10*/;
                       Tsco5_4_V_0 <= Tsi1_SPILL_257;
                       Tsin1_17_V_1 <= Tsi1_SPILL_257;
                       end 
                      
                  10'sd631/*631:xpc10*/:  begin 
                       xpc10 <= 10'sd208/*208:xpc10*/;
                       Tspr4_3_V_0 <= 64'sh8_0000_0000_0000|Tspr4_3_V_0;
                       end 
                      
                  10'sd632/*632:xpc10*/:  begin 
                       xpc10 <= 10'sd206/*206:xpc10*/;
                       Tspr4_3_V_3 <= (-64'sh20_0000_0000_0000<$signed((Tspr4_3_V_1<<32'sd1)));
                       end 
                      
                  10'sd634/*634:xpc10*/:  begin 
                       xpc10 <= 10'sd212/*212:xpc10*/;
                       Tsfl1_18_V_6 <= 64'shf_ffff_ffff_ffff&Tsf1_SPILL_256;
                       end 
                      
                  10'sd637/*637:xpc10*/:  begin 
                       xpc10 <= 10'sd638/*638:xpc10*/;
                       Tspr11_2_V_3 <= (-64'sh20_0000_0000_0000<$signed((Tspr11_2_V_1<<32'sd1)));
                       Tspr11_2_V_2 <= rtl_unsigned_bitextract5(Tsf0SPILL10_256);
                       end 
                      
                  10'sd639/*639:xpc10*/:  begin 
                       xpc10 <= 10'sd640/*640:xpc10*/;
                       Tspr11_2_V_0 <= 64'sh8_0000_0000_0000|Tspr11_2_V_0;
                       Tspr11_2_V_4 <= rtl_unsigned_bitextract5(Tsf0SPILL12_256);
                       end 
                      
                  10'sd640/*640:xpc10*/:  begin 
                       xpc10 <= 10'sd641/*641:xpc10*/;
                       Tspr11_2_V_1 <= 64'sh8_0000_0000_0000|Tspr11_2_V_1;
                       end 
                      
                  10'sd644/*644:xpc10*/:  begin 
                       xpc10 <= 10'sd640/*640:xpc10*/;
                       Tspr11_2_V_0 <= 64'sh8_0000_0000_0000|Tspr11_2_V_0;
                       end 
                      
                  10'sd645/*645:xpc10*/:  begin 
                       xpc10 <= 10'sd638/*638:xpc10*/;
                       Tspr11_2_V_3 <= (-64'sh20_0000_0000_0000<$signed((Tspr11_2_V_1<<32'sd1)));
                       end 
                      
                  10'sd652/*652:xpc10*/:  begin 
                       xpc10 <= 10'sd653/*653:xpc10*/;
                       Tsco3_7_V_0 <= (Tsco3_7_V_0<<32'sd8);
                       end 
                      
                  10'sd653/*653:xpc10*/:  begin 
                       xpc10 <= 10'sd654/*654:xpc10*/;
                       Tsco3_7_V_1 <= rtl_unsigned_bitextract3(Tsco3_7_V_1+A_8_US_CC_SCALbx14_ARA0[$unsigned((Tsco3_7_V_0>>32'sd24))]
                      );

                       end 
                      
                  10'sd654/*654:xpc10*/:  begin 
                       xpc10 <= 10'sd655/*655:xpc10*/;
                       Tsco0_2_V_1 <= rtl_unsigned_bitextract3(Tsco0_2_V_1+Tsco3_7_V_1);
                       end 
                      
                  10'sd655/*655:xpc10*/:  begin 
                       xpc10 <= 10'sd656/*656:xpc10*/;
                       Tsno19_4_V_0 <= $unsigned(-32'sd11+rtl_sign_extend10(Tsco0_2_V_1));
                       end 
                      
                  10'sd656/*656:xpc10*/:  begin 
                       xpc10 <= 10'sd657/*657:xpc10*/;
                       Tsfl1_7_V_6 <= (Tsfl1_7_V_6<<(32'sd63&Tsno19_4_V_0));
                       end 
                      
                  10'sd657/*657:xpc10*/:  begin 
                       xpc10 <= 10'sd658/*658:xpc10*/;
                       Tsfl1_7_V_3 <= rtl_signed_bitextract0(rtl_sign_extend2(16'sd1)+(0-Tsno19_4_V_0));
                       end 
                      
                  10'sd663/*663:xpc10*/:  begin 
                       xpc10 <= 10'sd664/*664:xpc10*/;
                       Tsco3_7_V_0 <= (Tsco3_7_V_0<<32'sd8);
                       end 
                      
                  10'sd664/*664:xpc10*/:  begin 
                       xpc10 <= 10'sd665/*665:xpc10*/;
                       Tsco3_7_V_1 <= rtl_unsigned_bitextract3(Tsco3_7_V_1+A_8_US_CC_SCALbx14_ARA0[$unsigned((Tsco3_7_V_0>>32'sd24))]
                      );

                       end 
                      
                  10'sd665/*665:xpc10*/:  begin 
                       xpc10 <= 10'sd666/*666:xpc10*/;
                       Tsco0_2_V_1 <= rtl_unsigned_bitextract3(Tsco0_2_V_1+Tsco3_7_V_1);
                       end 
                      
                  10'sd666/*666:xpc10*/:  begin 
                       xpc10 <= 10'sd667/*667:xpc10*/;
                       Tsno23_4_V_0 <= $unsigned(-32'sd11+rtl_sign_extend10(Tsco0_2_V_1));
                       end 
                      
                  10'sd667/*667:xpc10*/:  begin 
                       xpc10 <= 10'sd668/*668:xpc10*/;
                       Tsfl1_7_V_7 <= (Tsfl1_7_V_7<<(32'sd63&Tsno23_4_V_0));
                       end 
                      
                  10'sd668/*668:xpc10*/:  begin 
                       xpc10 <= 10'sd669/*669:xpc10*/;
                       Tsfl1_7_V_4 <= rtl_signed_bitextract0(rtl_sign_extend2(16'sd1)+(0-Tsno23_4_V_0));
                       end 
                      
                  10'sd669/*669:xpc10*/:  begin 
                       xpc10 <= 10'sd670/*670:xpc10*/;
                       Tsfl1_7_V_5 <= rtl_signed_bitextract0(-16'sd1023+Tsfl1_7_V_3+Tsfl1_7_V_4);
                       end 
                      
                  10'sd670/*670:xpc10*/:  begin 
                       xpc10 <= 10'sd671/*671:xpc10*/;
                       Tsfl1_7_V_6 <= ((64'sh10_0000_0000_0000|Tsfl1_7_V_6)<<32'sd10);
                       end 
                      
                  10'sd671/*671:xpc10*/:  begin 
                       xpc10 <= 10'sd672/*672:xpc10*/;
                       Tsfl1_7_V_7 <= ((64'sh10_0000_0000_0000|Tsfl1_7_V_7)<<32'sd11);
                       end 
                      
                  10'sd672/*672:xpc10*/:  begin 
                       xpc10 <= 10'sd673/*673:xpc10*/;
                       Tsmu24_24_V_1 <= rtl_unsigned_bitextract1(64'h_ffff_ffff&Tsfl1_7_V_6);
                       end 
                      
                  10'sd673/*673:xpc10*/:  begin 
                       xpc10 <= 10'sd674/*674:xpc10*/;
                       Tsmu24_24_V_0 <= rtl_unsigned_bitextract1((Tsfl1_7_V_6>>32'sd32));
                       end 
                      
                  10'sd674/*674:xpc10*/:  begin 
                       xpc10 <= 10'sd675/*675:xpc10*/;
                       Tsmu24_24_V_3 <= rtl_unsigned_bitextract1(64'h_ffff_ffff&Tsfl1_7_V_7);
                       end 
                      
                  10'sd675/*675:xpc10*/:  begin 
                       xpc10 <= 10'sd676/*676:xpc10*/;
                       Tsmu24_24_V_2 <= rtl_unsigned_bitextract1((Tsfl1_7_V_7>>32'sd32));
                       end 
                      
                  10'sd676/*676:xpc10*/:  begin 
                       xpc10 <= 10'sd677/*677:xpc10*/;
                       Tsmu24_24_V_7 <= rtl_unsigned_extend7(Tsmu24_24_V_1)*rtl_unsigned_extend7(Tsmu24_24_V_3);
                       end 
                      
                  10'sd677/*677:xpc10*/:  begin 
                       xpc10 <= 10'sd678/*678:xpc10*/;
                       Tsmu24_24_V_5 <= rtl_unsigned_extend7(Tsmu24_24_V_1)*rtl_unsigned_extend7(Tsmu24_24_V_2);
                       end 
                      
                  10'sd678/*678:xpc10*/:  begin 
                       xpc10 <= 10'sd679/*679:xpc10*/;
                       Tsmu24_24_V_6 <= rtl_unsigned_extend7(Tsmu24_24_V_0)*rtl_unsigned_extend7(Tsmu24_24_V_3);
                       end 
                      
                  10'sd679/*679:xpc10*/:  begin 
                       xpc10 <= 10'sd680/*680:xpc10*/;
                       Tsmu24_24_V_4 <= rtl_unsigned_extend7(Tsmu24_24_V_0)*rtl_unsigned_extend7(Tsmu24_24_V_2);
                       end 
                      
                  10'sd680/*680:xpc10*/:  begin 
                       xpc10 <= 10'sd681/*681:xpc10*/;
                       Tsmu24_24_V_5 <= Tsmu24_24_V_5+Tsmu24_24_V_6;
                       end 
                      
                  10'sd682/*682:xpc10*/:  begin 
                       xpc10 <= 10'sd683/*683:xpc10*/;
                       Tsm24_SPILL_264 <= Tsmu24_24_V_4;
                       fastspilldup26 <= Tsmu24_24_V_4;
                       end 
                      
                  10'sd684/*684:xpc10*/:  begin 
                       xpc10 <= 10'sd685/*685:xpc10*/;
                       Tsmu24_24_V_4 <= Tsm24_SPILL_257+(Tsm24_SPILL_259<<32'sd32)+(Tsmu24_24_V_5>>32'sd32);
                       end 
                      
                  10'sd685/*685:xpc10*/:  begin 
                       xpc10 <= 10'sd686/*686:xpc10*/;
                       Tsmu24_24_V_5 <= (Tsmu24_24_V_5<<32'sd32);
                       end 
                      
                  10'sd686/*686:xpc10*/:  begin 
                       xpc10 <= 10'sd687/*687:xpc10*/;
                       Tsmu24_24_V_7 <= Tsmu24_24_V_7+Tsmu24_24_V_5;
                       end 
                      
                  10'sd687/*687:xpc10*/:  begin 
                       xpc10 <= 10'sd688/*688:xpc10*/;
                       Tsm24_SPILL_263 <= Tsmu24_24_V_4;
                       fastspilldup28 <= Tsmu24_24_V_4;
                       end 
                      
                  10'sd689/*689:xpc10*/:  begin 
                       xpc10 <= 10'sd690/*690:xpc10*/;
                       Tsmu24_24_V_4 <= Tsm24_SPILL_260+Tsm24_SPILL_262;
                       end 
                      
                  10'sd690/*690:xpc10*/:  begin 
                       xpc10 <= 10'sd691/*691:xpc10*/;
                       Tsfl1_7_V_8 <= Tsmu24_24_V_4;
                       Tsfl1_7_V_9 <= Tsmu24_24_V_7;
                       end 
                      
                  10'sd691/*691:xpc10*/:  begin 
                       xpc10 <= 10'sd692/*692:xpc10*/;
                       Tsf1_SPILL_260 <= Tsfl1_7_V_8;
                       fastspilldup30 <= Tsfl1_7_V_8;
                       end 
                      
                  10'sd693/*693:xpc10*/:  begin 
                       xpc10 <= 10'sd694/*694:xpc10*/;
                       Tsfl1_7_V_8 <= Tsf1_SPILL_257|Tsf1_SPILL_259;
                       end 
                      
                  10'sd695/*695:xpc10*/:  begin 
                       xpc10 <= 10'sd696/*696:xpc10*/;
                       Tsfl1_7_V_5 <= rtl_signed_bitextract0(-16'sd1+Tsfl1_7_V_5);
                       end 
                      
                  10'sd696/*696:xpc10*/:  begin 
                       xpc10 <= 10'sd697/*697:xpc10*/;
                       Tsro29_4_V_1 <= Tsfl1_7_V_8;
                       Tsro29_4_V_0 <= rtl_signed_bitextract0(Tsfl1_7_V_5);
                       end 
                      
                  10'sd698/*698:xpc10*/:  begin 
                       xpc10 <= 10'sd699/*699:xpc10*/;
                       Tsro29_4_V_6 <= rtl_signed_bitextract9(64'sh3ff&Tsro29_4_V_1);
                       Tsro29_4_V_5 <= 16'sh200;
                       end 
                      
                  10'sd701/*701:xpc10*/:  begin 
                       xpc10 <= 10'sd702/*702:xpc10*/;
                       Tsr29_SPILL_256 <= fastspilldup32;
                       Tsr29_SPILL_260 <= fastspilldup32;
                       end 
                      
                  10'sd703/*703:xpc10*/:  begin 
                       xpc10 <= 10'sd704/*704:xpc10*/;
                       Tsr29_SPILL_259 <= Tsr29_SPILL_257+(0-Tsr29_SPILL_258);
                       end 
                      
                  10'sd705/*705:xpc10*/:  begin 
                       xpc10 <= 10'sd704/*704:xpc10*/;
                       Tsr29_SPILL_259 <= Tsr29_SPILL_257+(0-Tsr29_SPILL_258);
                       end 
                      
                  10'sd706/*706:xpc10*/:  begin 
                       xpc10 <= 10'sd707/*707:xpc10*/;
                       Tsro29_4_V_0 <= 16'sh0;
                       Tsro29_4_V_1 <= Tssh18_7_V_0;
                       end 
                      
                  10'sd707/*707:xpc10*/:  begin 
                       xpc10 <= 10'sd708/*708:xpc10*/;
                       Tsro29_4_V_6 <= rtl_signed_bitextract9(64'sh3ff&Tsro29_4_V_1);
                       end 
                      
                  10'sd710/*710:xpc10*/:  begin 
                       xpc10 <= 10'sd711/*711:xpc10*/;
                       Tsro29_4_V_1 <= (Tsro29_4_V_1+rtl_sign_extend4(Tsro29_4_V_5)>>32'sd10);
                       end 
                      
                  10'sd713/*713:xpc10*/:  begin 
                       xpc10 <= 10'sd714/*714:xpc10*/;
                       Tsr29_SPILL_259 <= Tsro29_4_V_1+(Tsp27_SPILL_256<<32'sd63)+(rtl_sign_extend4(Tsro29_4_V_0)<<32'sd52);
                       end 
                      
                  10'sd715/*715:xpc10*/:  begin 
                       xpc10 <= 10'sd714/*714:xpc10*/;
                       Tsr29_SPILL_259 <= Tsro29_4_V_1+(Tsp27_SPILL_256<<32'sd63)+(rtl_sign_extend4(Tsro29_4_V_0)<<32'sd52);
                       end 
                      
                  10'sd716/*716:xpc10*/:  begin 
                       xpc10 <= 10'sd717/*717:xpc10*/;
                       Tss18_SPILL_256 <= fastspilldup34;
                       Tss18_SPILL_259 <= fastspilldup34;
                       end 
                      
                  10'sd718/*718:xpc10*/:  begin 
                       xpc10 <= 10'sd719/*719:xpc10*/;
                       Tssh18_7_V_0 <= Tss18_SPILL_258|Tss18_SPILL_257;
                       end 
                      
                  10'sd719/*719:xpc10*/:  begin 
                       xpc10 <= 10'sd707/*707:xpc10*/;
                       Tsro29_4_V_0 <= 16'sh0;
                       Tsro29_4_V_1 <= Tssh18_7_V_0;
                       end 
                      
                  10'sd720/*720:xpc10*/:  begin 
                       xpc10 <= 10'sd719/*719:xpc10*/;
                       Tssh18_7_V_0 <= Tss18_SPILL_258|Tss18_SPILL_257;
                       end 
                      
                  10'sd721/*721:xpc10*/:  begin 
                       xpc10 <= 10'sd722/*722:xpc10*/;
                       Tsro29_4_V_1 <= Tss18_SPILL_260;
                       Tssh18_7_V_0 <= Tss18_SPILL_260;
                       end 
                      
                  10'sd722/*722:xpc10*/:  begin 
                       xpc10 <= 10'sd708/*708:xpc10*/;
                       Tsro29_4_V_6 <= rtl_signed_bitextract9(64'sh3ff&Tsro29_4_V_1);
                       Tsro29_4_V_0 <= 16'sh0;
                       end 
                      
                  10'sd723/*723:xpc10*/:  begin 
                       xpc10 <= 10'sd722/*722:xpc10*/;
                       Tsro29_4_V_1 <= Tss18_SPILL_260;
                       Tssh18_7_V_0 <= Tss18_SPILL_260;
                       end 
                      
                  10'sd724/*724:xpc10*/:  begin 
                       xpc10 <= 10'sd694/*694:xpc10*/;
                       Tsfl1_7_V_8 <= Tsf1_SPILL_260|Tsf1_SPILL_259;
                       end 
                      
                  10'sd725/*725:xpc10*/:  begin 
                       xpc10 <= 10'sd690/*690:xpc10*/;
                       Tsmu24_24_V_4 <= Tsm24_SPILL_263+Tsm24_SPILL_262;
                       end 
                      
                  10'sd726/*726:xpc10*/:  begin 
                       xpc10 <= 10'sd685/*685:xpc10*/;
                       Tsmu24_24_V_4 <= Tsm24_SPILL_264+(Tsm24_SPILL_259<<32'sd32)+(Tsmu24_24_V_5>>32'sd32);
                       end 
                      
                  10'sd727/*727:xpc10*/:  begin 
                       xpc10 <= 10'sd661/*661:xpc10*/;
                       Tsco3_7_V_0 <= rtl_unsigned_bitextract1(64'h_ffff_ffff&Tsco0_2_V_0);
                       end 
                      
                  10'sd728/*728:xpc10*/:  begin 
                       xpc10 <= 10'sd650/*650:xpc10*/;
                       Tsco3_7_V_0 <= rtl_unsigned_bitextract1(64'h_ffff_ffff&Tsco0_2_V_0);
                       end 
                      
                  10'sd729/*729:xpc10*/:  begin 
                       xpc10 <= 10'sd190/*190:xpc10*/;
                       Tspr4_3_V_0 <= 64'sh8_0000_0000_0000|Tspr4_3_V_0;
                       end 
                      
                  10'sd730/*730:xpc10*/:  begin 
                       xpc10 <= 10'sd188/*188:xpc10*/;
                       Tspr4_3_V_3 <= (-64'sh20_0000_0000_0000<$signed((Tspr4_3_V_1<<32'sd1)));
                       end 
                      
                  10'sd731/*731:xpc10*/:  begin 
                       xpc10 <= 10'sd194/*194:xpc10*/;
                       Tsfl0_10_V_0 <= 64'shff_ffff_ffff_ffff_ffff;
                       Tsf0_SPILL_256 <= 64'h_7fff_ffff_ffff_ffff;
                       end 
                      
                  10'sd732/*732:xpc10*/:  begin 
                       xpc10 <= 10'sd194/*194:xpc10*/;
                       Tsfl0_10_V_0 <= -64'sh_8000_0000_0000_0000&~Tsf0_SPILL_256|64'sh_7fff_ffff_ffff_ffff&Tsf0_SPILL_256;
                       end 
                      
                  10'sd733/*733:xpc10*/:  begin 
                       xpc10 <= 10'sd734/*734:xpc10*/;
                       Tspr11_2_V_1 <= $unsigned(A_64_US_CC_SCALbx12_ARB0[Tdbm0_3_V_1]);
                       end 
                      
                  10'sd735/*735:xpc10*/:  begin 
                       xpc10 <= 10'sd736/*736:xpc10*/;
                       Tspr11_2_V_3 <= (-64'sh20_0000_0000_0000<$signed((Tspr11_2_V_1<<32'sd1)));
                       Tspr11_2_V_2 <= rtl_unsigned_bitextract5(Tsf0SPILL10_256);
                       end 
                      
                  10'sd737/*737:xpc10*/:  begin 
                       xpc10 <= 10'sd738/*738:xpc10*/;
                       Tspr11_2_V_0 <= 64'sh8_0000_0000_0000|Tspr11_2_V_0;
                       Tspr11_2_V_4 <= rtl_unsigned_bitextract5(Tsf0SPILL12_256);
                       end 
                      
                  10'sd738/*738:xpc10*/:  begin 
                       xpc10 <= 10'sd739/*739:xpc10*/;
                       Tspr11_2_V_1 <= 64'sh8_0000_0000_0000|Tspr11_2_V_1;
                       end 
                      
                  10'sd741/*741:xpc10*/:  begin 
                       xpc10 <= 10'sd194/*194:xpc10*/;
                       Tsfl0_10_V_0 <= -64'sh_8000_0000_0000_0000&~Tsf0_SPILL_256|64'sh_7fff_ffff_ffff_ffff&Tsf0_SPILL_256;
                       end 
                      
                  10'sd742/*742:xpc10*/:  begin 
                       xpc10 <= 10'sd738/*738:xpc10*/;
                       Tspr11_2_V_0 <= 64'sh8_0000_0000_0000|Tspr11_2_V_0;
                       end 
                      
                  10'sd743/*743:xpc10*/:  begin 
                       xpc10 <= 10'sd736/*736:xpc10*/;
                       Tspr11_2_V_3 <= (-64'sh20_0000_0000_0000<$signed((Tspr11_2_V_1<<32'sd1)));
                       end 
                      
                  10'sd744/*744:xpc10*/:  begin 
                       xpc10 <= 10'sd194/*194:xpc10*/;
                       Tsfl0_10_V_0 <= 64'shff_ffff_ffff_ffff_ffff;
                       Tsf0_SPILL_256 <= 64'h_7fff_ffff_ffff_ffff;
                       end 
                      
                  10'sd745/*745:xpc10*/:  begin 
                       xpc10 <= 10'sd194/*194:xpc10*/;
                       Tsfl0_10_V_0 <= -64'sh_8000_0000_0000_0000&~Tsf0_SPILL_256|64'sh_7fff_ffff_ffff_ffff&Tsf0_SPILL_256;
                       end 
                      
                  10'sd746/*746:xpc10*/:  begin 
                       xpc10 <= 10'sd194/*194:xpc10*/;
                       Tsfl0_10_V_0 <= -64'sh_8000_0000_0000_0000&~Tsf0_SPILL_256|64'sh_7fff_ffff_ffff_ffff&Tsf0_SPILL_256;
                       end 
                      
                  10'sd750/*750:xpc10*/:  begin 
                       xpc10 <= 10'sd751/*751:xpc10*/;
                       Tsco3_7_V_0 <= (Tsco3_7_V_0<<32'sd8);
                       end 
                      
                  10'sd751/*751:xpc10*/:  begin 
                       xpc10 <= 10'sd752/*752:xpc10*/;
                       Tsco3_7_V_1 <= rtl_unsigned_bitextract3(Tsco3_7_V_1+A_8_US_CC_SCALbx14_ARA0[$unsigned((Tsco3_7_V_0>>32'sd24))]
                      );

                       end 
                      
                  10'sd752/*752:xpc10*/:  begin 
                       xpc10 <= 10'sd753/*753:xpc10*/;
                       Tsco0_2_V_1 <= rtl_unsigned_bitextract3(Tsco0_2_V_1+Tsco3_7_V_1);
                       end 
                      
                  10'sd753/*753:xpc10*/:  begin 
                       xpc10 <= 10'sd754/*754:xpc10*/;
                       Tsno19_4_V_0 <= $unsigned(-32'sd11+rtl_sign_extend10(Tsco0_2_V_1));
                       end 
                      
                  10'sd754/*754:xpc10*/:  begin 
                       xpc10 <= 10'sd755/*755:xpc10*/;
                       Tsfl0_9_V_6 <= (Tsfl0_9_V_6<<(32'sd63&Tsno19_4_V_0));
                       end 
                      
                  10'sd755/*755:xpc10*/:  begin 
                       xpc10 <= 10'sd756/*756:xpc10*/;
                       Tsfl0_9_V_3 <= rtl_signed_bitextract0(rtl_sign_extend2(16'sd1)+(0-Tsno19_4_V_0));
                       end 
                      
                  10'sd757/*757:xpc10*/:  begin 
                       xpc10 <= 10'sd194/*194:xpc10*/;
                       Tsfl0_10_V_0 <= -64'sh_8000_0000_0000_0000&~Tsf0_SPILL_256|64'sh_7fff_ffff_ffff_ffff&Tsf0_SPILL_256;
                       end 
                      
                  10'sd761/*761:xpc10*/:  begin 
                       xpc10 <= 10'sd762/*762:xpc10*/;
                       Tsco3_7_V_0 <= (Tsco3_7_V_0<<32'sd8);
                       end 
                      
                  10'sd762/*762:xpc10*/:  begin 
                       xpc10 <= 10'sd763/*763:xpc10*/;
                       Tsco3_7_V_1 <= rtl_unsigned_bitextract3(Tsco3_7_V_1+A_8_US_CC_SCALbx14_ARA0[$unsigned((Tsco3_7_V_0>>32'sd24))]
                      );

                       end 
                      
                  10'sd763/*763:xpc10*/:  begin 
                       xpc10 <= 10'sd764/*764:xpc10*/;
                       Tsco0_2_V_1 <= rtl_unsigned_bitextract3(Tsco0_2_V_1+Tsco3_7_V_1);
                       end 
                      
                  10'sd764/*764:xpc10*/:  begin 
                       xpc10 <= 10'sd765/*765:xpc10*/;
                       Tsno23_4_V_0 <= $unsigned(-32'sd11+rtl_sign_extend10(Tsco0_2_V_1));
                       end 
                      
                  10'sd765/*765:xpc10*/:  begin 
                       xpc10 <= 10'sd766/*766:xpc10*/;
                       Tsfl0_9_V_7 <= (Tsfl0_9_V_7<<(32'sd63&Tsno23_4_V_0));
                       end 
                      
                  10'sd766/*766:xpc10*/:  begin 
                       xpc10 <= 10'sd767/*767:xpc10*/;
                       Tsfl0_9_V_4 <= rtl_signed_bitextract0(rtl_sign_extend2(16'sd1)+(0-Tsno23_4_V_0));
                       end 
                      
                  10'sd767/*767:xpc10*/:  begin 
                       xpc10 <= 10'sd768/*768:xpc10*/;
                       Tsfl0_9_V_5 <= rtl_signed_bitextract0(-16'sd1023+Tsfl0_9_V_3+Tsfl0_9_V_4);
                       end 
                      
                  10'sd768/*768:xpc10*/:  begin 
                       xpc10 <= 10'sd769/*769:xpc10*/;
                       Tsfl0_9_V_6 <= ((64'sh10_0000_0000_0000|Tsfl0_9_V_6)<<32'sd10);
                       end 
                      
                  10'sd769/*769:xpc10*/:  begin 
                       xpc10 <= 10'sd770/*770:xpc10*/;
                       Tsfl0_9_V_7 <= ((64'sh10_0000_0000_0000|Tsfl0_9_V_7)<<32'sd11);
                       end 
                      
                  10'sd770/*770:xpc10*/:  begin 
                       xpc10 <= 10'sd771/*771:xpc10*/;
                       Tsmu24_24_V_1 <= rtl_unsigned_bitextract1(64'h_ffff_ffff&Tsfl0_9_V_6);
                       end 
                      
                  10'sd771/*771:xpc10*/:  begin 
                       xpc10 <= 10'sd772/*772:xpc10*/;
                       Tsmu24_24_V_0 <= rtl_unsigned_bitextract1((Tsfl0_9_V_6>>32'sd32));
                       end 
                      
                  10'sd772/*772:xpc10*/:  begin 
                       xpc10 <= 10'sd773/*773:xpc10*/;
                       Tsmu24_24_V_3 <= rtl_unsigned_bitextract1(64'h_ffff_ffff&Tsfl0_9_V_7);
                       end 
                      
                  10'sd773/*773:xpc10*/:  begin 
                       xpc10 <= 10'sd774/*774:xpc10*/;
                       Tsmu24_24_V_2 <= rtl_unsigned_bitextract1((Tsfl0_9_V_7>>32'sd32));
                       end 
                      
                  10'sd774/*774:xpc10*/:  begin 
                       xpc10 <= 10'sd775/*775:xpc10*/;
                       Tsmu24_24_V_7 <= rtl_unsigned_extend7(Tsmu24_24_V_1)*rtl_unsigned_extend7(Tsmu24_24_V_3);
                       end 
                      
                  10'sd775/*775:xpc10*/:  begin 
                       xpc10 <= 10'sd776/*776:xpc10*/;
                       Tsmu24_24_V_5 <= rtl_unsigned_extend7(Tsmu24_24_V_1)*rtl_unsigned_extend7(Tsmu24_24_V_2);
                       end 
                      
                  10'sd776/*776:xpc10*/:  begin 
                       xpc10 <= 10'sd777/*777:xpc10*/;
                       Tsmu24_24_V_6 <= rtl_unsigned_extend7(Tsmu24_24_V_0)*rtl_unsigned_extend7(Tsmu24_24_V_3);
                       end 
                      
                  10'sd777/*777:xpc10*/:  begin 
                       xpc10 <= 10'sd778/*778:xpc10*/;
                       Tsmu24_24_V_4 <= rtl_unsigned_extend7(Tsmu24_24_V_0)*rtl_unsigned_extend7(Tsmu24_24_V_2);
                       end 
                      
                  10'sd778/*778:xpc10*/:  begin 
                       xpc10 <= 10'sd779/*779:xpc10*/;
                       Tsmu24_24_V_5 <= Tsmu24_24_V_5+Tsmu24_24_V_6;
                       end 
                      
                  10'sd780/*780:xpc10*/:  begin 
                       xpc10 <= 10'sd781/*781:xpc10*/;
                       Tsm24_SPILL_264 <= Tsmu24_24_V_4;
                       fastspilldup16 <= Tsmu24_24_V_4;
                       end 
                      
                  10'sd782/*782:xpc10*/:  begin 
                       xpc10 <= 10'sd783/*783:xpc10*/;
                       Tsmu24_24_V_4 <= Tsm24_SPILL_257+(Tsm24_SPILL_259<<32'sd32)+(Tsmu24_24_V_5>>32'sd32);
                       end 
                      
                  10'sd783/*783:xpc10*/:  begin 
                       xpc10 <= 10'sd784/*784:xpc10*/;
                       Tsmu24_24_V_5 <= (Tsmu24_24_V_5<<32'sd32);
                       end 
                      
                  10'sd784/*784:xpc10*/:  begin 
                       xpc10 <= 10'sd785/*785:xpc10*/;
                       Tsmu24_24_V_7 <= Tsmu24_24_V_7+Tsmu24_24_V_5;
                       end 
                      
                  10'sd785/*785:xpc10*/:  begin 
                       xpc10 <= 10'sd786/*786:xpc10*/;
                       Tsm24_SPILL_263 <= Tsmu24_24_V_4;
                       fastspilldup18 <= Tsmu24_24_V_4;
                       end 
                      
                  10'sd787/*787:xpc10*/:  begin 
                       xpc10 <= 10'sd788/*788:xpc10*/;
                       Tsmu24_24_V_4 <= Tsm24_SPILL_260+Tsm24_SPILL_262;
                       end 
                      
                  10'sd788/*788:xpc10*/:  begin 
                       xpc10 <= 10'sd789/*789:xpc10*/;
                       Tsfl0_9_V_8 <= Tsmu24_24_V_4;
                       Tsfl0_9_V_9 <= Tsmu24_24_V_7;
                       end 
                      
                  10'sd789/*789:xpc10*/:  begin 
                       xpc10 <= 10'sd790/*790:xpc10*/;
                       Tsf0_SPILL_260 <= Tsfl0_9_V_8;
                       fastspilldup20 <= Tsfl0_9_V_8;
                       end 
                      
                  10'sd791/*791:xpc10*/:  begin 
                       xpc10 <= 10'sd792/*792:xpc10*/;
                       Tsfl0_9_V_8 <= Tsf0_SPILL_257|Tsf0_SPILL_259;
                       end 
                      
                  10'sd793/*793:xpc10*/:  begin 
                       xpc10 <= 10'sd794/*794:xpc10*/;
                       Tsfl0_9_V_5 <= rtl_signed_bitextract0(-16'sd1+Tsfl0_9_V_5);
                       end 
                      
                  10'sd794/*794:xpc10*/:  begin 
                       xpc10 <= 10'sd795/*795:xpc10*/;
                       Tsro29_4_V_1 <= Tsfl0_9_V_8;
                       Tsro29_4_V_0 <= rtl_signed_bitextract0(Tsfl0_9_V_5);
                       end 
                      
                  10'sd796/*796:xpc10*/:  begin 
                       xpc10 <= 10'sd797/*797:xpc10*/;
                       Tsro29_4_V_6 <= rtl_signed_bitextract9(64'sh3ff&Tsro29_4_V_1);
                       Tsro29_4_V_5 <= 16'sh200;
                       end 
                      
                  10'sd799/*799:xpc10*/:  begin 
                       xpc10 <= 10'sd800/*800:xpc10*/;
                       Tsr29_SPILL_256 <= fastspilldup22;
                       Tsr29_SPILL_260 <= fastspilldup22;
                       end 
                      
                  10'sd801/*801:xpc10*/:  begin 
                       xpc10 <= 10'sd802/*802:xpc10*/;
                       Tsr29_SPILL_259 <= Tsr29_SPILL_257+(0-Tsr29_SPILL_258);
                       end 
                      
                  10'sd802/*802:xpc10*/:  begin 
                       xpc10 <= 10'sd194/*194:xpc10*/;
                       Tsfl0_10_V_0 <= -64'sh_8000_0000_0000_0000&~Tsr29_SPILL_259|64'sh_7fff_ffff_ffff_ffff&Tsr29_SPILL_259;
                       Tsf0_SPILL_256 <= Tsr29_SPILL_259;
                       end 
                      
                  10'sd803/*803:xpc10*/:  begin 
                       xpc10 <= 10'sd802/*802:xpc10*/;
                       Tsr29_SPILL_259 <= Tsr29_SPILL_257+(0-Tsr29_SPILL_258);
                       end 
                      
                  10'sd804/*804:xpc10*/:  begin 
                       xpc10 <= 10'sd805/*805:xpc10*/;
                       Tsro29_4_V_0 <= 16'sh0;
                       Tsro29_4_V_1 <= Tssh18_7_V_0;
                       end 
                      
                  10'sd805/*805:xpc10*/:  begin 
                       xpc10 <= 10'sd806/*806:xpc10*/;
                       Tsro29_4_V_6 <= rtl_signed_bitextract9(64'sh3ff&Tsro29_4_V_1);
                       end 
                      
                  10'sd808/*808:xpc10*/:  begin 
                       xpc10 <= 10'sd809/*809:xpc10*/;
                       Tsro29_4_V_1 <= (Tsro29_4_V_1+rtl_sign_extend4(Tsro29_4_V_5)>>32'sd10);
                       end 
                      
                  10'sd811/*811:xpc10*/:  begin 
                       xpc10 <= 10'sd812/*812:xpc10*/;
                       Tsr29_SPILL_259 <= Tsro29_4_V_1+(Tsp27_SPILL_256<<32'sd63)+(rtl_sign_extend4(Tsro29_4_V_0)<<32'sd52);
                       end 
                      
                  10'sd812/*812:xpc10*/:  begin 
                       xpc10 <= 10'sd194/*194:xpc10*/;
                       Tsfl0_10_V_0 <= -64'sh_8000_0000_0000_0000&~Tsr29_SPILL_259|64'sh_7fff_ffff_ffff_ffff&Tsr29_SPILL_259;
                       Tsf0_SPILL_256 <= Tsr29_SPILL_259;
                       end 
                      
                  10'sd813/*813:xpc10*/:  begin 
                       xpc10 <= 10'sd812/*812:xpc10*/;
                       Tsr29_SPILL_259 <= Tsro29_4_V_1+(Tsp27_SPILL_256<<32'sd63)+(rtl_sign_extend4(Tsro29_4_V_0)<<32'sd52);
                       end 
                      
                  10'sd814/*814:xpc10*/:  begin 
                       xpc10 <= 10'sd815/*815:xpc10*/;
                       Tss18_SPILL_256 <= fastspilldup24;
                       Tss18_SPILL_259 <= fastspilldup24;
                       end 
                      
                  10'sd816/*816:xpc10*/:  begin 
                       xpc10 <= 10'sd817/*817:xpc10*/;
                       Tssh18_7_V_0 <= Tss18_SPILL_258|Tss18_SPILL_257;
                       end 
                      
                  10'sd817/*817:xpc10*/:  begin 
                       xpc10 <= 10'sd805/*805:xpc10*/;
                       Tsro29_4_V_0 <= 16'sh0;
                       Tsro29_4_V_1 <= Tssh18_7_V_0;
                       end 
                      
                  10'sd818/*818:xpc10*/:  begin 
                       xpc10 <= 10'sd817/*817:xpc10*/;
                       Tssh18_7_V_0 <= Tss18_SPILL_258|Tss18_SPILL_257;
                       end 
                      
                  10'sd819/*819:xpc10*/:  begin 
                       xpc10 <= 10'sd820/*820:xpc10*/;
                       Tsro29_4_V_1 <= Tss18_SPILL_260;
                       Tssh18_7_V_0 <= Tss18_SPILL_260;
                       end 
                      
                  10'sd820/*820:xpc10*/:  begin 
                       xpc10 <= 10'sd806/*806:xpc10*/;
                       Tsro29_4_V_6 <= rtl_signed_bitextract9(64'sh3ff&Tsro29_4_V_1);
                       Tsro29_4_V_0 <= 16'sh0;
                       end 
                      
                  10'sd821/*821:xpc10*/:  begin 
                       xpc10 <= 10'sd820/*820:xpc10*/;
                       Tsro29_4_V_1 <= Tss18_SPILL_260;
                       Tssh18_7_V_0 <= Tss18_SPILL_260;
                       end 
                      
                  10'sd822/*822:xpc10*/:  begin 
                       xpc10 <= 10'sd792/*792:xpc10*/;
                       Tsfl0_9_V_8 <= Tsf0_SPILL_260|Tsf0_SPILL_259;
                       end 
                      
                  10'sd823/*823:xpc10*/:  begin 
                       xpc10 <= 10'sd788/*788:xpc10*/;
                       Tsmu24_24_V_4 <= Tsm24_SPILL_263+Tsm24_SPILL_262;
                       end 
                      
                  10'sd824/*824:xpc10*/:  begin 
                       xpc10 <= 10'sd783/*783:xpc10*/;
                       Tsmu24_24_V_4 <= Tsm24_SPILL_264+(Tsm24_SPILL_259<<32'sd32)+(Tsmu24_24_V_5>>32'sd32);
                       end 
                      
                  10'sd825/*825:xpc10*/:  begin 
                       xpc10 <= 10'sd759/*759:xpc10*/;
                       Tsco3_7_V_0 <= rtl_unsigned_bitextract1(64'h_ffff_ffff&Tsco0_2_V_0);
                       end 
                      
                  10'sd826/*826:xpc10*/:  begin 
                       xpc10 <= 10'sd748/*748:xpc10*/;
                       Tsco3_7_V_0 <= rtl_unsigned_bitextract1(64'h_ffff_ffff&Tsco0_2_V_0);
                       end 
                      endcase
              if ((xpc10==10'sd20/*20:xpc10*/))  xpc10 <= 10'sd21/*21:xpc10*/;
                  if ((xpc10==10'sd40/*40:xpc10*/))  xpc10 <= 10'sd41/*41:xpc10*/;
                  if ((xpc10==10'sd170/*170:xpc10*/))  xpc10 <= 10'sd171/*171:xpc10*/;
                  if ((xpc10==10'sd173/*173:xpc10*/))  xpc10 <= 10'sd174/*174:xpc10*/;
                  if ((xpc10==10'sd274/*274:xpc10*/))  xpc10 <= 10'sd275/*275:xpc10*/;
                  if ((xpc10==10'sd378/*378:xpc10*/))  xpc10 <= 10'sd379/*379:xpc10*/;
                  if ((xpc10==10'sd517/*517:xpc10*/))  xpc10 <= 10'sd518/*518:xpc10*/;
                  if ((xpc10==10'sd536/*536:xpc10*/))  xpc10 <= 10'sd537/*537:xpc10*/;
                  if ((xpc10==10'sd584/*584:xpc10*/))  xpc10 <= 10'sd585/*585:xpc10*/;
                  if ((xpc10==10'sd681/*681:xpc10*/))  xpc10 <= 10'sd682/*682:xpc10*/;
                  if ((xpc10==10'sd697/*697:xpc10*/))  xpc10 <= 10'sd698/*698:xpc10*/;
                  if ((xpc10==10'sd779/*779:xpc10*/))  xpc10 <= 10'sd780/*780:xpc10*/;
                  if ((xpc10==10'sd795/*795:xpc10*/))  xpc10 <= 10'sd796/*796:xpc10*/;
                   end 
              //End structure HPR dfsin


       end 
      

// 1 vectors of width 10
// 207 vectors of width 64
// 48 vectors of width 1
// 27 vectors of width 16
// 15 vectors of width 32
// 3 vectors of width 8
// 72 array locations of width 64
// 259 array locations of width 8
// 768 bits in scalar variables
// Total state bits in module = 21690 bits.
// Total number of leaf cells = 0
endmodule

//  
// LCP delay estimations included: turn off with -vnl-lcp-delay-estimate=disable
//HPR L/S (orangepath) auxiliary reports.
//KiwiC compilation report
//Kiwi Scientific Acceleration (KiwiC .net/CIL/C# to Verilog/SystemC compiler): Version alpha 0.2.16f : 22nd-September-2016
//25/09/2016 22:35:42
//Cmd line args:  /home/djg11/d320/hprls/kiwipro/kiwic/distro/lib/kiwic.exe -vnl-resets=synchronous -restructure2=disable -vnl-roundtrip=disable -kiwic-cil-dump=combined -kiwic-kcode-dump=enable -bevelab-default-pause-mode=soft -bevelab-soft-pause-threshold=10 dfsin.exe -vnl=dfsin.v -vnl-resets=synchronous ../softfloat.dll


//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation KiKiwi for prefix KiwiSystem/Kiwi

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation SyBitConverter for prefix System/BitConverter

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation CS0.4 for prefix CS/0.4

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation @8 for prefix @/8

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation CS0.10 for prefix CS/0.10

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation @64 for prefix @/64

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tdb0._SPILL for prefix T404/dfsin/bm_main/0.3/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tdbm0.3 for prefix T404/dfsin/bm_main/0.3

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tdsi3.5 for prefix T404/dfsin/sin/3.5

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsf0._SPILL for prefix T404/softfloat/float64_mul/0.9/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsfl0.9 for prefix T404/softfloat/float64_mul/0.9

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tse0._SPILL for prefix T404/softfloat/extractFloat64Sign/0.14/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tse0SPILL10 for prefix T404/softfloat/extractFloat64Sign/0.23/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsp4._SPILL for prefix T404/softfloat/propagateFloat64NaN/4.3/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tspr4.3 for prefix T404/softfloat/propagateFloat64NaN/4.3

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsf0SPILL10 for prefix T404/softfloat/float64_is_signaling_nan/0.6/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsf0SPILL12 for prefix T404/softfloat/float64_is_signaling_nan/0.12/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsp8._SPILL for prefix T404/softfloat/packFloat64/8.5/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsp11_SPILL for prefix T404/softfloat/propagateFloat64NaN/11.2/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tspr11.2 for prefix T404/softfloat/propagateFloat64NaN/11.2

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsp15_SPILL for prefix T404/softfloat/packFloat64/15.5/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsp18_SPILL for prefix T404/softfloat/packFloat64/18.4/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsno19.4 for prefix T404/softfloat/normalizeFloat64Subnormal/19.4

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsco0.2 for prefix T404/softfloat/countLeadingZeros64/0.2

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsco3.7 for prefix T404/softfloat/countLeadingZeros32/3.7

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsp22_SPILL for prefix T404/softfloat/packFloat64/22.4/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsno23.4 for prefix T404/softfloat/normalizeFloat64Subnormal/23.4

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsm24_SPILL for prefix T404/softfloat/mul64To128/24.24/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsmu24.24 for prefix T404/softfloat/mul64To128/24.24

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsr29_SPILL for prefix T404/softfloat/roundAndPackFloat64/29.4/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsro29.4 for prefix T404/softfloat/roundAndPackFloat64/29.4

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsp13_SPILL for prefix T404/softfloat/packFloat64/13.7/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tss18_SPILL for prefix T404/softfloat/shift64RightJamming/18.7/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tssh18.7 for prefix T404/softfloat/shift64RightJamming/18.7

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsp27_SPILL for prefix T404/softfloat/packFloat64/27.4/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsfl0.10 for prefix T404/softfloat/float64_neg/0.10

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsf1._SPILL for prefix T404/softfloat/float64_mul/1.7/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsfl1.7 for prefix T404/softfloat/float64_mul/1.7

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsi1._SPILL for prefix T404/softfloat/int32_to_float64/1.17/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsin1.17 for prefix T404/softfloat/int32_to_float64/1.17

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsco5.4 for prefix T404/softfloat/countLeadingZeros32/5.4

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsp5._SPILL for prefix T404/softfloat/packFloat64/5.21/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsf1SPILL10 for prefix T404/softfloat/float64_div/1.18/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsfl1.18 for prefix T404/softfloat/float64_div/1.18

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tse0SPILL12 for prefix T404/softfloat/extractFloat64Sign/0.8/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tse0SPILL14 for prefix T404/softfloat/extractFloat64Sign/0.17/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsp2._SPILL for prefix T404/softfloat/propagateFloat64NaN/2.2/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tspr2.2 for prefix T404/softfloat/propagateFloat64NaN/2.2

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsp5SPILL10 for prefix T404/softfloat/propagateFloat64NaN/5.2/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tspr5.2 for prefix T404/softfloat/propagateFloat64NaN/5.2

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsp7._SPILL for prefix T404/softfloat/packFloat64/7.5/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsp10_SPILL for prefix T404/softfloat/propagateFloat64NaN/10.2/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tspr10.2 for prefix T404/softfloat/propagateFloat64NaN/10.2

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsp11SPILL10 for prefix T404/softfloat/packFloat64/11.5/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsp17_SPILL for prefix T404/softfloat/packFloat64/17.7/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsno18.4 for prefix T404/softfloat/normalizeFloat64Subnormal/18.4

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsp21_SPILL for prefix T404/softfloat/packFloat64/21.4/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsno22.4 for prefix T404/softfloat/normalizeFloat64Subnormal/22.4

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tse25_SPILL for prefix T404/softfloat/estimateDiv128To64/25.5/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tses25.5 for prefix T404/softfloat/estimateDiv128To64/25.5

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsm5._SPILL for prefix T404/softfloat/mul64To128/5.7/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsmu5.7 for prefix T404/softfloat/mul64To128/5.7

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tss5._SPILL for prefix T404/softfloat/sub128/5.14/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsa6._SPILL for prefix T404/softfloat/add128/6.15/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsad6.15 for prefix T404/softfloat/add128/6.15

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsm26_SPILL for prefix T404/softfloat/mul64To128/26.4/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsmu26.4 for prefix T404/softfloat/mul64To128/26.4

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tss26_SPILL for prefix T404/softfloat/sub128/26.12/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsa27_SPILL for prefix T404/softfloat/add128/27.13/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsad27.13 for prefix T404/softfloat/add128/27.13

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsr33_SPILL for prefix T404/softfloat/roundAndPackFloat64/33.4/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsro33.4 for prefix T404/softfloat/roundAndPackFloat64/33.4

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsf1SPILL12 for prefix T404/softfloat/float64_add/1.22/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsfl1.22 for prefix T404/softfloat/float64_add/1.22

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tse0SPILL16 for prefix T404/softfloat/extractFloat64Sign/0.2/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tse0SPILL18 for prefix T404/softfloat/extractFloat64Sign/0.5/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsa1._SPILL for prefix T404/softfloat/addFloat64Sigs/1.3/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsad1.3 for prefix T404/softfloat/addFloat64Sigs/1.3

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsp3._SPILL for prefix T404/softfloat/propagateFloat64NaN/3.2/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tspr3.2 for prefix T404/softfloat/propagateFloat64NaN/3.2

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tss8._SPILL for prefix T404/softfloat/shift64RightJamming/8.5/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tssh8.5 for prefix T404/softfloat/shift64RightJamming/8.5

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsp12_SPILL for prefix T404/softfloat/propagateFloat64NaN/12.2/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tspr12.2 for prefix T404/softfloat/propagateFloat64NaN/12.2

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsp13SPILL10 for prefix T404/softfloat/packFloat64/13.5/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tss17_SPILL for prefix T404/softfloat/shift64RightJamming/17.6/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tssh17.6 for prefix T404/softfloat/shift64RightJamming/17.6

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsp21SPILL10 for prefix T404/softfloat/propagateFloat64NaN/21.3/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tspr21.3 for prefix T404/softfloat/propagateFloat64NaN/21.3

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsp24_SPILL for prefix T404/softfloat/packFloat64/24.7/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsr28_SPILL for prefix T404/softfloat/roundAndPackFloat64/28.4/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsro28.4 for prefix T404/softfloat/roundAndPackFloat64/28.4

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tss2._SPILL for prefix T404/softfloat/subFloat64Sigs/2.4/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tssu2.4 for prefix T404/softfloat/subFloat64Sigs/2.4

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsp7SPILL10 for prefix T404/softfloat/propagateFloat64NaN/7.3/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tspr7.3 for prefix T404/softfloat/propagateFloat64NaN/7.3

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsp18SPILL10 for prefix T404/softfloat/propagateFloat64NaN/18.2/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tspr18.2 for prefix T404/softfloat/propagateFloat64NaN/18.2

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsp19_SPILL for prefix T404/softfloat/packFloat64/19.7/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tss23_SPILL for prefix T404/softfloat/shift64RightJamming/23.6/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tssh23.6 for prefix T404/softfloat/shift64RightJamming/23.6

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsp27SPILL10 for prefix T404/softfloat/propagateFloat64NaN/27.2/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tspr27.2 for prefix T404/softfloat/propagateFloat64NaN/27.2

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tss32_SPILL for prefix T404/softfloat/shift64RightJamming/32.5/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tssh32.5 for prefix T404/softfloat/shift64RightJamming/32.5

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsno34.9 for prefix T404/softfloat/normalizeRoundAndPackFloat64/34.9

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsr0._SPILL for prefix T404/softfloat/roundAndPackFloat64/0.16/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsro0.16 for prefix T404/softfloat/roundAndPackFloat64/0.16

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsf0SPILL14 for prefix T404/softfloat/float64_le/0.3/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsfl0.3 for prefix T404/softfloat/float64_le/0.3

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tse5._SPILL for prefix T404/softfloat/extractFloat64Sign/5.2/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tse5SPILL10 for prefix T404/softfloat/extractFloat64Sign/5.5/_SPILL

//----------------------------------------------------------

//Report from KiwiC-fe.rpt:::
//KiwiC: front end input processing of class or method called KiwiSystem/Kiwi
//
//root_walk start thread at a static method (used as an entry point). Method name=.cctor uid=cctor10
//
//KiwiC start_thread (or entry point) id=cctor10
//
//Root method elaborated: specificf=S_kickoff_collate leftover=1+0
//
//KiwiC: front end input processing of class or method called System/BitConverter
//
//root_walk start thread at a static method (used as an entry point). Method name=.cctor uid=cctor12
//
//KiwiC start_thread (or entry point) id=cctor12
//
//Root method elaborated: specificf=S_kickoff_collate leftover=1+1
//
//KiwiC: front end input processing of class or method called softfloat
//
//root_walk start thread at a static method (used as an entry point). Method name=.cctor uid=cctor14
//
//KiwiC start_thread (or entry point) id=cctor14
//
//Root method elaborated: specificf=S_kickoff_collate leftover=1+2
//
//KiwiC: front end input processing of class or method called dfsin
//
//root_walk start thread at a static method (used as an entry point). Method name=.cctor uid=cctor16
//
//KiwiC start_thread (or entry point) id=cctor16
//
//Root method elaborated: specificf=S_kickoff_collate leftover=1+3
//
//KiwiC: front end input processing of class or method called dfsin
//
//root_compiler: start elaborating class 'dfsin'
//
//elaborating class 'dfsin'
//
//compiling static method as entry point: style=Root idl=dfsin/HWMain
//
//Performing root elaboration of method HWMain
//
//KiwiC start_thread (or entry point) id=HWMain10
//
//root_compiler class done: dfsin
//
//Report of all settings used from the recipe or command line:
//
//   cil-uwind-budget=10000
//
//   kiwic-finish=enable
//
//   kiwic-cil-dump=combined
//
//   kiwic-kcode-dump=enable
//
//   kiwic-register-colours=disable
//
//   array-4d-name=KIWIARRAY4D
//
//   array-3d-name=KIWIARRAY3D
//
//   array-2d-name=KIWIARRAY2D
//
//   kiwi-dll=Kiwi.dll
//
//   kiwic-dll=Kiwic.dll
//
//   kiwic-zerolength-arrays=disable
//
//   kiwic-fpgaconsole-default=enable
//
//   postgen-optimise=enable
//
//   gtrace-loglevel=20
//
//   firstpass-loglevel=20
//
//   root=$attributeroot
//
//   ?>?=srcfile, dfsin.exe, ../softfloat.dll
//
//END OF KIWIC REPORT FILE
//

//----------------------------------------------------------

//Report from enumbers:::
//Concise expression alias report.
//
//  -- No expression aliases to report
//

//----------------------------------------------------------

//Report from verilog_render:::
//1 vectors of width 10
//
//207 vectors of width 64
//
//48 vectors of width 1
//
//27 vectors of width 16
//
//15 vectors of width 32
//
//3 vectors of width 8
//
//72 array locations of width 64
//
//259 array locations of width 8
//
//768 bits in scalar variables
//
//Total state bits in module = 21690 bits.
//
//Total number of leaf cells = 0
//

//Major Statistics Report:
//Thread .cctor uid=cctor10 has 3 CIL instructions in 1 basic blocks
//Thread .cctor uid=cctor12 has 2 CIL instructions in 1 basic blocks
//Thread .cctor uid=cctor14 has 6 CIL instructions in 1 basic blocks
//Thread .cctor uid=cctor16 has 11 CIL instructions in 1 basic blocks
//Thread HWMain uid=HWMain10 has 2201 CIL instructions in 851 basic blocks
//Thread mpc10 has 827 bevelab control states (pauses)
// eof (HPR L/S Verilog)
