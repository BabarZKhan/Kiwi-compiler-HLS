

// CBG Orangepath HPR L/S System

// Verilog output file generated at 30/03/2016 09:24:20
// Kiwi Scientific Acceleration (KiwiC .net/CIL/C# to Verilog/SystemC compiler): Version alpha 2.06: 22-Mar-2016 Unix 3.19.8.100
//  /home/djg11/d320/hprls/kiwipro/kiwic/distro/lib/kiwic.exe -vnl-roundtrip=disable -report-each-step -kiwic-finish=enable -kiwic-kcode-dump=enable test44.exe -sim 1800 -vnl-resets=synchronous -vnl test44.v -res2-no-dram-ports=0 -give-backtrace -report-each-step
`timescale 1ns/10ps


module test44(input clk, input reset);
// Total state bits in module = 0 bits.
// Total number of leaf cells = 0
endmodule

// 
/*

// Restructure Technology Settings
*------------------------+---------+---------------------------------------------------------------------------------*
| Key                    | Value   | Description                                                                     |
*------------------------+---------+---------------------------------------------------------------------------------*
| int_flr_mul            | 16000   |                                                                                 |
| fp_fl_dp_div           | 5       |                                                                                 |
| fp_fl_dp_add           | 5       |                                                                                 |
| fp_fl_dp_mul           | 5       |                                                                                 |
| fp_fl_sp_div           | 5       |                                                                                 |
| fp_fl_sp_add           | 5       |                                                                                 |
| fp_fl_sp_mul           | 5       |                                                                                 |
| max_no_fp_muls         | 6       | Maximum number of adders and subtractors (or combos) to instantiate per thread. |
| max_no_fp_muls         | 6       | Maximum number of f/p dividers to instantiate per thread.                       |
| max_no_int_muls        | 3       | Maximum number of int multipliers to instantiate per thread.                    |
| max_no_fp_divs         | 2       | Maximum number of f/p dividers to instantiate per thread.                       |
| max_no_int_divs        | 2       | Maximum number of int dividers to instantiate per thread.                       |
| res2-offchip-threshold | 1000000 |                                                                                 |
| res2-combram-threshold | 32      |                                                                                 |
| res2-regfile-threshold | 8       |                                                                                 |
*------------------------+---------+---------------------------------------------------------------------------------*

// Offchip Memory Physical Ports/Banks = Nothing to Report

// */

//  
// LCP delay estimations included: turn off with -vnl-lcp-delay-estimate=disable
// eof (HPR L/S Verilog)
