

// CBG Orangepath HPR L/S System

// Verilog output file generated at 23/09/2016 20:09:06
// Kiwi Scientific Acceleration (KiwiC .net/CIL/C# to Verilog/SystemC compiler): Version alpha 0.2.16f : 22nd-September-2016 Linux/X86_64:koo
//  /home/djg11/d320/hprls/kiwipro/kiwic/distro/lib/kiwic.exe -vnl-resets=synchronous -restructure2=disable -vnl-roundtrip=disable -kiwic-cil-dump=combined -kiwic-kcode-dump=enable -bevelab-default-pause-mode=maximal -bevelab-soft-pause-threshold=10 dfsin.exe ../softfloat.dll
`timescale 1ns/1ns


module dfsin(output reg done, input [31:0] dfsin_arg, output [31:0] dfsin_result, input clk, input reset);
function signed [15:0] rtl_signed_bitextract2;
   input [63:0] arg;
   rtl_signed_bitextract2 = $signed(arg[15:0]);
   endfunction

function signed [15:0] rtl_signed_bitextract0;
   input [31:0] arg;
   rtl_signed_bitextract0 = $signed(arg[15:0]);
   endfunction

function  rtl_unsigned_bitextract12;
   input [31:0] arg;
   rtl_unsigned_bitextract12 = $unsigned(arg[0:0]);
   endfunction

function [7:0] rtl_unsigned_bitextract7;
   input [31:0] arg;
   rtl_unsigned_bitextract7 = $unsigned(arg[7:0]);
   endfunction

function [31:0] rtl_unsigned_bitextract6;
   input [63:0] arg;
   rtl_unsigned_bitextract6 = $unsigned(arg[31:0]);
   endfunction

function  rtl_unsigned_bitextract4;
   input [31:0] arg;
   rtl_unsigned_bitextract4 = $unsigned(arg[0:0]);
   endfunction

function signed [63:0] rtl_sign_extend11;
   input [15:0] arg;
   rtl_sign_extend11 = { {48{arg[15]}}, arg[15:0] };
   endfunction

function signed [31:0] rtl_sign_extend9;
   input [15:0] arg;
   rtl_sign_extend9 = { {16{arg[15]}}, arg[15:0] };
   endfunction

function signed [31:0] rtl_sign_extend8;
   input [7:0] arg;
   rtl_sign_extend8 = { {24{arg[7]}}, arg[7:0] };
   endfunction

function signed [63:0] rtl_sign_extend5;
   input argbit;
   rtl_sign_extend5 = { {64{argbit}} };
   endfunction

function signed [31:0] rtl_sign_extend3;
   input argbit;
   rtl_sign_extend3 = { {32{argbit}} };
   endfunction

function signed [63:0] rtl_sign_extend1;
   input [31:0] arg;
   rtl_sign_extend1 = { {32{arg[31]}}, arg[31:0] };
   endfunction

function [63:0] rtl_unsigned_extend10;
   input [31:0] arg;
   rtl_unsigned_extend10 = { 32'b0, arg[31:0] };
   endfunction

  integer Tdbm0_3_V_0;
  integer Tdbm0_3_V_1;
  reg [63:0] Tdsi1_5_V_0;
  reg [63:0] Tdsi1_5_V_1;
  integer Tdsi1_5_V_2;
  reg [63:0] Tsfl0_9_V_8;
  reg [63:0] Tsfl0_9_V_9;
  reg [63:0] Tsfl0_9_V_6;
  reg signed [15:0] Tsfl0_9_V_3;
  integer Tse0_SPILL_256;
  reg Tsfl0_9_V_0;
  reg [63:0] Tsfl0_9_V_7;
  reg signed [15:0] Tsfl0_9_V_4;
  integer Tse0SPILL10_256;
  reg Tsfl0_9_V_1;
  reg Tsfl0_9_V_2;
  reg [63:0] Tsf0_SPILL_256;
  reg signed [63:0] Tsp8_SPILL_256;
  reg [63:0] Tspr4_3_V_0;
  reg [63:0] Tspr4_3_V_1;
  integer Tsf0SPILL10_256;
  reg Tspr4_3_V_2;
  reg Tspr4_3_V_3;
  integer Tsf0SPILL12_256;
  reg Tspr4_3_V_4;
  reg [63:0] Tsp4_SPILL_256;
  reg [63:0] Tspr11_2_V_0;
  reg [63:0] Tspr11_2_V_1;
  reg Tspr11_2_V_2;
  reg Tspr11_2_V_3;
  reg Tspr11_2_V_4;
  reg [63:0] Tsp11_SPILL_256;
  reg signed [63:0] Tsp15_SPILL_256;
  reg signed [63:0] Tsp18_SPILL_256;
  reg [63:0] Tsco0_2_V_0;
  reg [7:0] Tsco0_2_V_1;
  reg [31:0] Tsco3_7_V_0;
  reg [7:0] Tsco3_7_V_1;
  integer Tsno19_4_V_0;
  reg signed [63:0] Tsp22_SPILL_256;
  integer Tsno23_4_V_0;
  reg signed [15:0] Tsfl0_9_V_5;
  reg [31:0] Tsmu24_24_V_1;
  reg [31:0] Tsmu24_24_V_0;
  reg [31:0] Tsmu24_24_V_3;
  reg [31:0] Tsmu24_24_V_2;
  reg [63:0] Tsmu24_24_V_7;
  reg [63:0] Tsmu24_24_V_5;
  reg [63:0] Tsmu24_24_V_6;
  reg [63:0] Tsmu24_24_V_4;
  reg [63:0] fastspilldup18;
  reg [63:0] Tsm24_SPILL_264;
  reg [63:0] Tsm24_SPILL_257;
  reg signed [63:0] Tsm24_SPILL_259;
  reg [63:0] Tsm24_SPILL_258;
  reg [63:0] fastspilldup20;
  reg [63:0] Tsm24_SPILL_263;
  reg [63:0] Tsm24_SPILL_260;
  reg signed [63:0] Tsm24_SPILL_262;
  reg [63:0] Tsm24_SPILL_261;
  reg [63:0] fastspilldup22;
  reg [63:0] Tsf0_SPILL_260;
  reg [63:0] Tsf0_SPILL_257;
  reg signed [63:0] Tsf0_SPILL_259;
  reg [63:0] Tsf0_SPILL_258;
  reg signed [15:0] Tsro29_4_V_0;
  reg [63:0] Tsro29_4_V_1;
  reg signed [15:0] Tsro29_4_V_5;
  reg signed [15:0] Tsro29_4_V_6;
  reg [63:0] Tssh18_7_V_0;
  reg [63:0] fastspilldup26;
  reg [63:0] Tss18_SPILL_259;
  reg [63:0] Tss18_SPILL_256;
  reg signed [63:0] Tss18_SPILL_258;
  reg [63:0] Tss18_SPILL_257;
  reg signed [63:0] Tss18_SPILL_260;
  reg signed [63:0] Tsp13_SPILL_256;
  reg [63:0] fastspilldup24;
  reg [63:0] Tsr29_SPILL_260;
  reg [63:0] Tsr29_SPILL_256;
  reg signed [63:0] Tsr29_SPILL_258;
  reg [63:0] Tsr29_SPILL_257;
  reg [63:0] Tsr29_SPILL_259;
  reg signed [63:0] Tsp27_SPILL_256;
  reg [63:0] Tsfl0_10_V_0;
  reg [63:0] Tdsi1_5_V_3;
  reg [63:0] Tsfl1_8_V_8;
  reg [63:0] Tsfl1_8_V_9;
  reg [63:0] Tsfl1_8_V_6;
  reg signed [15:0] Tsfl1_8_V_3;
  reg Tsfl1_8_V_0;
  reg [63:0] Tsfl1_8_V_7;
  reg signed [15:0] Tsfl1_8_V_4;
  reg Tsfl1_8_V_1;
  reg Tsfl1_8_V_2;
  reg [63:0] Tsf1_SPILL_256;
  reg signed [15:0] Tsfl1_8_V_5;
  reg [63:0] fastspilldup28;
  reg [63:0] fastspilldup30;
  reg [63:0] fastspilldup32;
  reg [63:0] Tsf1_SPILL_260;
  reg [63:0] Tsf1_SPILL_257;
  reg signed [63:0] Tsf1_SPILL_259;
  reg [63:0] Tsf1_SPILL_258;
  reg [63:0] fastspilldup36;
  reg [63:0] fastspilldup34;
  reg [63:0] Tsi1_SPILL_256;
  reg Tsin1_19_V_0;
  integer Tsi1_SPILL_257;
  reg [31:0] Tsin1_19_V_1;
  reg [31:0] Tsco5_4_V_0;
  reg [7:0] Tsco5_4_V_1;
  integer Tsin1_19_V_3;
  reg [63:0] Tsin1_19_V_2;
  reg signed [63:0] Tsp5_SPILL_256;
  reg [63:0] Tsfl1_24_V_8;
  reg [63:0] Tsfl1_24_V_9;
  reg [63:0] Tsfl1_24_V_6;
  reg signed [15:0] Tsfl1_24_V_3;
  reg Tsfl1_24_V_0;
  reg [63:0] Tsfl1_24_V_7;
  reg signed [15:0] Tsfl1_24_V_4;
  reg Tsfl1_24_V_1;
  reg Tsfl1_24_V_2;
  reg [63:0] Tsf1SPILL10_256;
  reg signed [15:0] Tsfl1_24_V_5;
  reg [63:0] fastspilldup38;
  reg [63:0] fastspilldup40;
  reg [63:0] fastspilldup42;
  reg [63:0] Tsf1SPILL10_260;
  reg [63:0] Tsf1SPILL10_257;
  reg signed [63:0] Tsf1SPILL10_259;
  reg [63:0] Tsf1SPILL10_258;
  reg [63:0] fastspilldup46;
  reg [63:0] fastspilldup44;
  reg [63:0] Tsi1SPILL10_256;
  reg Tsin1_34_V_0;
  integer Tsi1SPILL10_257;
  reg [31:0] Tsin1_34_V_1;
  integer Tsin1_34_V_3;
  reg [63:0] Tsin1_34_V_2;
  reg [63:0] Tsfl1_35_V_6;
  reg signed [15:0] Tsfl1_35_V_3;
  integer Tse0SPILL12_256;
  reg Tsfl1_35_V_0;
  reg [63:0] Tsfl1_35_V_7;
  reg signed [15:0] Tsfl1_35_V_4;
  integer Tse0SPILL14_256;
  reg Tsfl1_35_V_1;
  reg Tsfl1_35_V_2;
  reg [63:0] Tspr2_2_V_0;
  reg [63:0] Tspr2_2_V_1;
  reg Tspr2_2_V_2;
  reg Tspr2_2_V_3;
  reg Tspr2_2_V_4;
  reg [63:0] Tsp2_SPILL_256;
  reg [63:0] Tsf1SPILL12_256;
  reg [63:0] Tspr5_2_V_0;
  reg [63:0] Tspr5_2_V_1;
  reg Tspr5_2_V_2;
  reg Tspr5_2_V_3;
  reg Tspr5_2_V_4;
  reg [63:0] Tsp5SPILL10_256;
  reg signed [63:0] Tsp7_SPILL_256;
  reg [63:0] Tspr10_2_V_0;
  reg [63:0] Tspr10_2_V_1;
  reg Tspr10_2_V_2;
  reg Tspr10_2_V_3;
  reg Tspr10_2_V_4;
  reg [63:0] Tsp10_SPILL_256;
  reg signed [63:0] Tsp11SPILL10_256;
  reg signed [63:0] Tsp17_SPILL_256;
  integer Tsno18_4_V_0;
  reg signed [63:0] Tsp21_SPILL_256;
  integer Tsno22_4_V_0;
  reg signed [15:0] Tsfl1_35_V_5;
  reg [63:0] Tse25_SPILL_256;
  reg [63:0] Tses25_5_V_0;
  reg [63:0] Tse25_SPILL_257;
  reg [63:0] Tses25_5_V_6;
  reg [31:0] Tsmu5_7_V_1;
  reg [31:0] Tsmu5_7_V_0;
  reg [31:0] Tsmu5_7_V_3;
  reg [31:0] Tsmu5_7_V_2;
  reg [63:0] Tsmu5_7_V_7;
  reg [63:0] Tsmu5_7_V_5;
  reg [63:0] Tsmu5_7_V_6;
  reg [63:0] Tsmu5_7_V_4;
  reg [63:0] fastspilldup48;
  reg [63:0] Tsm5_SPILL_264;
  reg [63:0] Tsm5_SPILL_257;
  reg signed [63:0] Tsm5_SPILL_259;
  reg [63:0] Tsm5_SPILL_258;
  reg [63:0] fastspilldup50;
  reg [63:0] Tsm5_SPILL_263;
  reg [63:0] Tsm5_SPILL_260;
  reg signed [63:0] Tsm5_SPILL_262;
  reg [63:0] Tsm5_SPILL_261;
  reg [63:0] Tses25_5_V_5;
  reg [63:0] Tses25_5_V_4;
  reg [63:0] Tses25_5_V_3;
  reg [63:0] fastspilldup52;
  reg [63:0] Tss5_SPILL_262;
  reg [63:0] Tss5_SPILL_257;
  reg signed [63:0] Tss5_SPILL_260;
  reg [63:0] Tss5_SPILL_259;
  reg [63:0] Tses25_5_V_2;
  reg [63:0] fastspilldup56;
  reg [63:0] Tse25_SPILL_261;
  reg [63:0] Tse25_SPILL_258;
  reg [63:0] Tse25_SPILL_260;
  reg [63:0] Tse25_SPILL_259;
  reg [63:0] Tsfl1_35_V_8;
  reg [31:0] Tsmu26_4_V_1;
  reg [31:0] Tsmu26_4_V_0;
  reg [31:0] Tsmu26_4_V_3;
  reg [31:0] Tsmu26_4_V_2;
  reg [63:0] Tsmu26_4_V_7;
  reg [63:0] Tsmu26_4_V_5;
  reg [63:0] Tsmu26_4_V_6;
  reg [63:0] Tsmu26_4_V_4;
  reg [63:0] fastspilldup58;
  reg [63:0] Tsm26_SPILL_264;
  reg [63:0] Tsm26_SPILL_257;
  reg signed [63:0] Tsm26_SPILL_259;
  reg [63:0] Tsm26_SPILL_258;
  reg [63:0] fastspilldup60;
  reg [63:0] Tsm26_SPILL_263;
  reg [63:0] Tsm26_SPILL_260;
  reg signed [63:0] Tsm26_SPILL_262;
  reg [63:0] Tsm26_SPILL_261;
  reg [63:0] Tsfl1_35_V_12;
  reg [63:0] Tsfl1_35_V_11;
  reg [63:0] Tsfl1_35_V_10;
  reg [63:0] fastspilldup62;
  reg [63:0] Tss26_SPILL_262;
  reg [63:0] Tss26_SPILL_257;
  reg signed [63:0] Tss26_SPILL_260;
  reg [63:0] Tss26_SPILL_259;
  reg [63:0] Tsfl1_35_V_9;
  reg [63:0] fastspilldup66;
  reg [63:0] Tsf1SPILL12_260;
  reg [63:0] Tsf1SPILL12_257;
  reg signed [63:0] Tsf1SPILL12_259;
  reg [63:0] Tsf1SPILL12_258;
  reg [63:0] Tsad27_13_V_0;
  reg [63:0] fastspilldup64;
  reg [63:0] Tsa27_SPILL_262;
  reg [63:0] Tsa27_SPILL_257;
  reg signed [63:0] Tsa27_SPILL_260;
  reg [63:0] Tsa27_SPILL_259;
  reg signed [15:0] Tsro33_4_V_0;
  reg [63:0] Tsro33_4_V_1;
  reg signed [15:0] Tsro33_4_V_5;
  reg signed [15:0] Tsro33_4_V_6;
  reg [63:0] fastspilldup70;
  reg [63:0] fastspilldup68;
  reg [63:0] Tsr33_SPILL_260;
  reg [63:0] Tsr33_SPILL_256;
  reg signed [63:0] Tsr33_SPILL_258;
  reg [63:0] Tsr33_SPILL_257;
  reg [63:0] Tsr33_SPILL_259;
  integer Tse0SPILL16_256;
  reg Tsfl1_39_V_0;
  integer Tse0SPILL18_256;
  reg Tsfl1_39_V_1;
  reg [63:0] Tsad1_3_V_3;
  reg signed [15:0] Tsad1_3_V_0;
  reg [63:0] Tsad1_3_V_4;
  reg signed [15:0] Tsad1_3_V_1;
  integer Tsad1_3_V_6;
  reg [63:0] Tspr3_2_V_0;
  reg [63:0] Tspr3_2_V_1;
  reg Tspr3_2_V_2;
  reg Tspr3_2_V_3;
  reg Tspr3_2_V_4;
  reg [63:0] Tsp3_SPILL_256;
  reg [63:0] Tsa1_SPILL_256;
  reg [63:0] Tssh8_5_V_0;
  reg [63:0] fastspilldup72;
  reg [63:0] Tss8_SPILL_259;
  reg [63:0] Tss8_SPILL_256;
  reg signed [63:0] Tss8_SPILL_258;
  reg [63:0] Tss8_SPILL_257;
  reg signed [63:0] Tss8_SPILL_260;
  reg signed [15:0] Tsad1_3_V_2;
  reg [63:0] Tspr12_2_V_0;
  reg [63:0] Tspr12_2_V_1;
  reg Tspr12_2_V_2;
  reg Tspr12_2_V_3;
  reg Tspr12_2_V_4;
  reg [63:0] Tsp12_SPILL_256;
  reg signed [63:0] Tsp13SPILL10_256;
  reg [63:0] Tssh17_6_V_0;
  reg [63:0] fastspilldup74;
  reg [63:0] Tss17_SPILL_259;
  reg [63:0] Tss17_SPILL_256;
  reg signed [63:0] Tss17_SPILL_258;
  reg [63:0] Tss17_SPILL_257;
  reg signed [63:0] Tss17_SPILL_260;
  reg [63:0] Tsad1_3_V_5;
  reg [63:0] Tspr21_3_V_0;
  reg [63:0] Tspr21_3_V_1;
  reg Tspr21_3_V_2;
  reg Tspr21_3_V_3;
  reg Tspr21_3_V_4;
  reg [63:0] Tsp21SPILL10_256;
  reg signed [63:0] Tsp24_SPILL_256;
  reg signed [15:0] Tsro28_4_V_0;
  reg [63:0] Tsro28_4_V_1;
  reg signed [15:0] Tsro28_4_V_5;
  reg signed [15:0] Tsro28_4_V_6;
  reg [63:0] fastspilldup78;
  reg [63:0] fastspilldup76;
  reg [63:0] Tsr28_SPILL_260;
  reg [63:0] Tsr28_SPILL_256;
  reg signed [63:0] Tsr28_SPILL_258;
  reg [63:0] Tsr28_SPILL_257;
  reg [63:0] Tsr28_SPILL_259;
  reg [63:0] Tsf1SPILL14_256;
  reg Tssu2_4_V_0;
  reg [63:0] Tssu2_4_V_4;
  reg signed [15:0] Tssu2_4_V_1;
  reg [63:0] Tssu2_4_V_5;
  reg signed [15:0] Tssu2_4_V_2;
  integer Tssu2_4_V_7;
  reg [63:0] Tspr27_2_V_0;
  reg [63:0] Tspr27_2_V_1;
  reg Tspr27_2_V_2;
  reg Tspr27_2_V_3;
  reg Tspr27_2_V_4;
  reg [63:0] Tsp27SPILL10_256;
  reg [63:0] Tss2_SPILL_256;
  reg [63:0] Tssh32_5_V_0;
  reg [63:0] fastspilldup82;
  reg [63:0] Tss32_SPILL_259;
  reg [63:0] Tss32_SPILL_256;
  reg signed [63:0] Tss32_SPILL_258;
  reg [63:0] Tss32_SPILL_257;
  reg signed [63:0] Tss32_SPILL_260;
  reg [63:0] Tspr18_2_V_0;
  reg [63:0] Tspr18_2_V_1;
  reg Tspr18_2_V_2;
  reg Tspr18_2_V_3;
  reg Tspr18_2_V_4;
  reg [63:0] Tsp18SPILL10_256;
  reg signed [63:0] Tsp19_SPILL_256;
  reg [63:0] Tssh23_6_V_0;
  reg [63:0] fastspilldup80;
  reg [63:0] Tss23_SPILL_259;
  reg [63:0] Tss23_SPILL_256;
  reg signed [63:0] Tss23_SPILL_258;
  reg [63:0] Tss23_SPILL_257;
  reg signed [63:0] Tss23_SPILL_260;
  reg [63:0] Tspr7_3_V_0;
  reg [63:0] Tspr7_3_V_1;
  reg Tspr7_3_V_2;
  reg Tspr7_3_V_3;
  reg Tspr7_3_V_4;
  reg [63:0] Tsp7SPILL10_256;
  reg [63:0] Tssu2_4_V_6;
  reg signed [15:0] Tssu2_4_V_3;
  integer Tsno34_9_V_0;
  reg signed [15:0] Tsro0_16_V_0;
  reg [63:0] Tsro0_16_V_1;
  reg signed [15:0] Tsro0_16_V_5;
  reg signed [15:0] Tsro0_16_V_6;
  reg [63:0] fastspilldup86;
  reg [63:0] fastspilldup84;
  reg [63:0] Tsr0_SPILL_260;
  reg [63:0] Tsr0_SPILL_256;
  reg signed [63:0] Tsr0_SPILL_258;
  reg [63:0] Tsr0_SPILL_257;
  reg [63:0] Tsr0_SPILL_259;
  integer Tsf0SPILL14_256;
  integer Tse5_SPILL_256;
  reg Tsfl0_3_V_0;
  integer Tse5SPILL10_256;
  reg Tsfl0_3_V_1;
  integer Tsf0SPILL14_257;
  integer Tsf0SPILL14_258;
  reg [63:0] Tdbm0_3_V_2;
  integer fastspilldup88;
  integer Tdb0_SPILL_259;
  integer Tdb0_SPILL_256;
  integer Tdb0_SPILL_258;
  integer Tdb0_SPILL_257;
  reg [63:0] Tses25_5_V_1;
  reg [63:0] Tsad6_15_V_0;
  reg [63:0] fastspilldup54;
  reg [63:0] Tsa6_SPILL_262;
  reg [63:0] Tsa6_SPILL_257;
  reg signed [63:0] Tsa6_SPILL_260;
  reg [63:0] Tsa6_SPILL_259;
  reg [7:0] A_8_US_CC_SCALbx16_ARA0[258:0];
  reg [63:0] A_64_US_CC_SCALbx12_ARB0[35:0];
  reg [63:0] A_64_US_CC_SCALbx10_ARA0[35:0];
  reg [12:0] xpc10;
 always   @(posedge clk )  begin 
      //Start structure HPR dfsin
      if (reset)  begin 
               Tsfl0_9_V_0 <= 32'd0;
               Tsfl0_9_V_1 <= 32'd0;
               Tsfl0_9_V_2 <= 32'd0;
               Tsfl0_10_V_0 <= 64'd0;
               Tdsi1_5_V_3 <= 64'd0;
               Tsfl1_8_V_0 <= 32'd0;
               Tsfl1_8_V_1 <= 32'd0;
               Tsfl1_8_V_2 <= 32'd0;
               Tsfl1_24_V_0 <= 32'd0;
               Tsfl1_24_V_1 <= 32'd0;
               Tsfl1_24_V_2 <= 32'd0;
               Tspr4_3_V_2 <= 32'd0;
               Tspr4_3_V_3 <= 32'd0;
               Tspr4_3_V_4 <= 32'd0;
               Tspr4_3_V_0 <= 64'd0;
               Tspr4_3_V_1 <= 64'd0;
               Tsfl1_35_V_0 <= 32'd0;
               Tsfl1_35_V_1 <= 32'd0;
               Tsfl1_35_V_2 <= 32'd0;
               Tspr2_2_V_2 <= 32'd0;
               Tspr2_2_V_3 <= 32'd0;
               Tspr2_2_V_4 <= 32'd0;
               Tspr2_2_V_0 <= 64'd0;
               Tspr2_2_V_1 <= 64'd0;
               Tdsi1_5_V_1 <= 64'd0;
               Tsfl1_39_V_0 <= 32'd0;
               Tsfl1_39_V_1 <= 32'd0;
               Tsad1_3_V_0 <= 32'd0;
               Tsad1_3_V_1 <= 32'd0;
               Tspr3_2_V_2 <= 32'd0;
               Tspr3_2_V_3 <= 32'd0;
               Tspr3_2_V_4 <= 32'd0;
               Tspr3_2_V_0 <= 64'd0;
               Tspr3_2_V_1 <= 64'd0;
               Tdsi1_5_V_0 <= 64'd0;
               Tdsi1_5_V_2 <= 32'd0;
               Tdbm0_3_V_2 <= 64'd0;
               fastspilldup88 <= 32'd0;
               Tdb0_SPILL_259 <= 32'd0;
               Tdb0_SPILL_256 <= 32'd0;
               Tdbm0_3_V_0 <= 32'd0;
               Tdbm0_3_V_1 <= 32'd0;
               done <= 32'd0;
               Tdb0_SPILL_258 <= 32'd0;
               Tdb0_SPILL_257 <= 32'd0;
               Tse5_SPILL_256 <= 32'd0;
               Tsfl0_3_V_0 <= 32'd0;
               Tsfl0_3_V_1 <= 32'd0;
               Tsf0SPILL14_257 <= 32'd0;
               Tsf0SPILL14_256 <= 32'd0;
               Tsf0SPILL14_258 <= 32'd0;
               Tse5SPILL10_256 <= 32'd0;
               Tsp3_SPILL_256 <= 64'd0;
               Tsro28_4_V_5 <= 32'd0;
               fastspilldup76 <= 64'd0;
               Tsr28_SPILL_260 <= 64'd0;
               Tsr28_SPILL_256 <= 64'd0;
               Tsr28_SPILL_258 <= 64'd0;
               Tsr28_SPILL_257 <= 64'd0;
               Tsro28_4_V_6 <= 32'd0;
               Tsro28_4_V_1 <= 64'd0;
               Tsro28_4_V_0 <= 32'd0;
               Tsr28_SPILL_259 <= 64'd0;
               fastspilldup78 <= 64'd0;
               fastspilldup72 <= 64'd0;
               Tss8_SPILL_259 <= 64'd0;
               Tss8_SPILL_256 <= 64'd0;
               Tss8_SPILL_258 <= 64'd0;
               Tss8_SPILL_257 <= 64'd0;
               Tssh8_5_V_0 <= 64'd0;
               Tss8_SPILL_260 <= 64'd0;
               Tsad1_3_V_4 <= 64'd0;
               Tspr12_2_V_2 <= 32'd0;
               Tspr12_2_V_3 <= 32'd0;
               Tspr12_2_V_4 <= 32'd0;
               Tspr12_2_V_0 <= 64'd0;
               Tspr12_2_V_1 <= 64'd0;
               Tsp12_SPILL_256 <= 64'd0;
               Tsp13SPILL10_256 <= 64'd0;
               Tsad1_3_V_6 <= 32'd0;
               fastspilldup74 <= 64'd0;
               Tss17_SPILL_259 <= 64'd0;
               Tss17_SPILL_256 <= 64'd0;
               Tss17_SPILL_258 <= 64'd0;
               Tss17_SPILL_257 <= 64'd0;
               Tssh17_6_V_0 <= 64'd0;
               Tss17_SPILL_260 <= 64'd0;
               Tsad1_3_V_3 <= 64'd0;
               Tspr21_3_V_2 <= 32'd0;
               Tspr21_3_V_3 <= 32'd0;
               Tspr21_3_V_4 <= 32'd0;
               Tspr21_3_V_0 <= 64'd0;
               Tspr21_3_V_1 <= 64'd0;
               Tsp21SPILL10_256 <= 64'd0;
               Tsa1_SPILL_256 <= 64'd0;
               Tsp24_SPILL_256 <= 64'd0;
               Tsad1_3_V_5 <= 64'd0;
               Tsad1_3_V_2 <= 32'd0;
               Tspr27_2_V_2 <= 32'd0;
               Tspr27_2_V_3 <= 32'd0;
               Tspr27_2_V_4 <= 32'd0;
               Tspr27_2_V_0 <= 64'd0;
               Tspr27_2_V_1 <= 64'd0;
               Tsf1SPILL14_256 <= 64'd0;
               Tsp27SPILL10_256 <= 64'd0;
               Tsno34_9_V_0 <= 32'd0;
               Tsro0_16_V_5 <= 32'd0;
               fastspilldup84 <= 64'd0;
               Tsr0_SPILL_260 <= 64'd0;
               Tsr0_SPILL_256 <= 64'd0;
               Tsr0_SPILL_258 <= 64'd0;
               Tsr0_SPILL_257 <= 64'd0;
               Tsro0_16_V_6 <= 32'd0;
               Tsro0_16_V_1 <= 64'd0;
               Tsro0_16_V_0 <= 32'd0;
               Tsr0_SPILL_259 <= 64'd0;
               fastspilldup86 <= 64'd0;
               fastspilldup82 <= 64'd0;
               Tss32_SPILL_259 <= 64'd0;
               Tss32_SPILL_256 <= 64'd0;
               Tss32_SPILL_258 <= 64'd0;
               Tss32_SPILL_257 <= 64'd0;
               Tssh32_5_V_0 <= 64'd0;
               Tss32_SPILL_260 <= 64'd0;
               Tspr18_2_V_2 <= 32'd0;
               Tspr18_2_V_3 <= 32'd0;
               Tspr18_2_V_4 <= 32'd0;
               Tspr18_2_V_0 <= 64'd0;
               Tspr18_2_V_1 <= 64'd0;
               Tsp18SPILL10_256 <= 64'd0;
               Tsp19_SPILL_256 <= 64'd0;
               Tssu2_4_V_7 <= 32'd0;
               Tssu2_4_V_5 <= 64'd0;
               Tssu2_4_V_6 <= 64'd0;
               Tssu2_4_V_3 <= 32'd0;
               Tssu2_4_V_0 <= 32'd0;
               fastspilldup80 <= 64'd0;
               Tss23_SPILL_259 <= 64'd0;
               Tss23_SPILL_256 <= 64'd0;
               Tss23_SPILL_258 <= 64'd0;
               Tss23_SPILL_257 <= 64'd0;
               Tssh23_6_V_0 <= 64'd0;
               Tss23_SPILL_260 <= 64'd0;
               Tssu2_4_V_4 <= 64'd0;
               Tspr7_3_V_2 <= 32'd0;
               Tspr7_3_V_3 <= 32'd0;
               Tspr7_3_V_4 <= 32'd0;
               Tspr7_3_V_0 <= 64'd0;
               Tspr7_3_V_1 <= 64'd0;
               Tsp7SPILL10_256 <= 64'd0;
               Tssu2_4_V_1 <= 32'd0;
               Tssu2_4_V_2 <= 32'd0;
               Tss2_SPILL_256 <= 64'd0;
               Tse0SPILL18_256 <= 32'd0;
               Tse0SPILL16_256 <= 32'd0;
               Tsp2_SPILL_256 <= 64'd0;
               Tspr5_2_V_2 <= 32'd0;
               Tspr5_2_V_3 <= 32'd0;
               Tspr5_2_V_4 <= 32'd0;
               Tspr5_2_V_0 <= 64'd0;
               Tspr5_2_V_1 <= 64'd0;
               Tsp5SPILL10_256 <= 64'd0;
               Tsp7_SPILL_256 <= 64'd0;
               Tspr10_2_V_2 <= 32'd0;
               Tspr10_2_V_3 <= 32'd0;
               Tspr10_2_V_4 <= 32'd0;
               Tspr10_2_V_0 <= 64'd0;
               Tspr10_2_V_1 <= 64'd0;
               Tsp10_SPILL_256 <= 64'd0;
               Tsp11SPILL10_256 <= 64'd0;
               Tsp17_SPILL_256 <= 64'd0;
               Tsno18_4_V_0 <= 32'd0;
               Tsfl1_35_V_4 <= 32'd0;
               Tsp21_SPILL_256 <= 64'd0;
               Tsno22_4_V_0 <= 32'd0;
               Tsfl1_35_V_3 <= 32'd0;
               Tsfl1_35_V_7 <= 64'd0;
               Tsfl1_35_V_6 <= 64'd0;
               Tsfl1_35_V_5 <= 32'd0;
               Tsmu26_4_V_1 <= 32'd0;
               Tsmu26_4_V_0 <= 32'd0;
               Tsmu26_4_V_3 <= 32'd0;
               Tsmu26_4_V_2 <= 32'd0;
               Tsmu26_4_V_6 <= 64'd0;
               fastspilldup58 <= 64'd0;
               Tsm26_SPILL_264 <= 64'd0;
               Tsm26_SPILL_257 <= 64'd0;
               Tsmu26_4_V_5 <= 64'd0;
               Tsmu26_4_V_7 <= 64'd0;
               fastspilldup60 <= 64'd0;
               Tsm26_SPILL_263 <= 64'd0;
               Tsm26_SPILL_260 <= 64'd0;
               Tsmu26_4_V_4 <= 64'd0;
               Tsfl1_35_V_12 <= 64'd0;
               Tsfl1_35_V_11 <= 64'd0;
               fastspilldup62 <= 64'd0;
               Tss26_SPILL_262 <= 64'd0;
               Tss26_SPILL_257 <= 64'd0;
               fastspilldup66 <= 64'd0;
               Tsf1SPILL12_260 <= 64'd0;
               Tsf1SPILL12_257 <= 64'd0;
               Tsro33_4_V_5 <= 32'd0;
               fastspilldup68 <= 64'd0;
               Tsr33_SPILL_260 <= 64'd0;
               Tsr33_SPILL_256 <= 64'd0;
               Tsf1SPILL12_256 <= 64'd0;
               Tsr33_SPILL_258 <= 64'd0;
               Tsr33_SPILL_257 <= 64'd0;
               Tsro33_4_V_6 <= 32'd0;
               Tsro33_4_V_1 <= 64'd0;
               Tsro33_4_V_0 <= 32'd0;
               Tsr33_SPILL_259 <= 64'd0;
               fastspilldup70 <= 64'd0;
               Tsf1SPILL12_259 <= 64'd0;
               Tsf1SPILL12_258 <= 64'd0;
               Tsfl1_35_V_8 <= 64'd0;
               Tsad27_13_V_0 <= 64'd0;
               Tsfl1_35_V_10 <= 64'd0;
               fastspilldup64 <= 64'd0;
               Tsa27_SPILL_262 <= 64'd0;
               Tsa27_SPILL_257 <= 64'd0;
               Tsfl1_35_V_9 <= 64'd0;
               Tsa27_SPILL_260 <= 64'd0;
               Tsa27_SPILL_259 <= 64'd0;
               Tss26_SPILL_260 <= 64'd0;
               Tss26_SPILL_259 <= 64'd0;
               Tsm26_SPILL_262 <= 64'd0;
               Tsm26_SPILL_261 <= 64'd0;
               Tsm26_SPILL_259 <= 64'd0;
               Tsm26_SPILL_258 <= 64'd0;
               Tses25_5_V_0 <= 64'd0;
               Tsmu5_7_V_1 <= 32'd0;
               Tsmu5_7_V_0 <= 32'd0;
               Tsmu5_7_V_3 <= 32'd0;
               Tsmu5_7_V_2 <= 32'd0;
               Tsmu5_7_V_6 <= 64'd0;
               fastspilldup48 <= 64'd0;
               Tsm5_SPILL_264 <= 64'd0;
               Tsm5_SPILL_257 <= 64'd0;
               Tsmu5_7_V_5 <= 64'd0;
               Tsmu5_7_V_7 <= 64'd0;
               fastspilldup50 <= 64'd0;
               Tsm5_SPILL_263 <= 64'd0;
               Tsm5_SPILL_260 <= 64'd0;
               Tsmu5_7_V_4 <= 64'd0;
               Tses25_5_V_5 <= 64'd0;
               Tses25_5_V_4 <= 64'd0;
               fastspilldup52 <= 64'd0;
               Tss5_SPILL_262 <= 64'd0;
               Tss5_SPILL_257 <= 64'd0;
               fastspilldup56 <= 64'd0;
               Tse25_SPILL_261 <= 64'd0;
               Tse25_SPILL_258 <= 64'd0;
               Tse25_SPILL_256 <= 64'd0;
               Tse25_SPILL_260 <= 64'd0;
               Tse25_SPILL_259 <= 64'd0;
               Tses25_5_V_6 <= 64'd0;
               Tses25_5_V_1 <= 64'd0;
               Tsad6_15_V_0 <= 64'd0;
               Tses25_5_V_3 <= 64'd0;
               fastspilldup54 <= 64'd0;
               Tsa6_SPILL_262 <= 64'd0;
               Tsa6_SPILL_257 <= 64'd0;
               Tses25_5_V_2 <= 64'd0;
               Tsa6_SPILL_260 <= 64'd0;
               Tsa6_SPILL_259 <= 64'd0;
               Tss5_SPILL_260 <= 64'd0;
               Tss5_SPILL_259 <= 64'd0;
               Tsm5_SPILL_262 <= 64'd0;
               Tsm5_SPILL_261 <= 64'd0;
               Tsm5_SPILL_259 <= 64'd0;
               Tsm5_SPILL_258 <= 64'd0;
               Tse25_SPILL_257 <= 64'd0;
               Tse0SPILL14_256 <= 32'd0;
               Tse0SPILL12_256 <= 32'd0;
               Tsin1_34_V_0 <= 32'd0;
               Tsin1_34_V_1 <= 32'd0;
               Tsin1_34_V_3 <= 32'd0;
               Tsin1_34_V_2 <= 64'd0;
               Tsi1SPILL10_256 <= 64'd0;
               Tsi1SPILL10_257 <= 32'd0;
               Tsfl1_24_V_3 <= 32'd0;
               Tsfl1_24_V_4 <= 32'd0;
               Tsfl1_24_V_6 <= 64'd0;
               Tsfl1_24_V_7 <= 64'd0;
               fastspilldup38 <= 64'd0;
               fastspilldup40 <= 64'd0;
               Tsfl1_24_V_9 <= 64'd0;
               fastspilldup42 <= 64'd0;
               Tsf1SPILL10_260 <= 64'd0;
               Tsf1SPILL10_257 <= 64'd0;
               Tsfl1_24_V_8 <= 64'd0;
               Tsfl1_24_V_5 <= 32'd0;
               fastspilldup44 <= 64'd0;
               Tsf1SPILL10_256 <= 64'd0;
               fastspilldup46 <= 64'd0;
               Tsf1SPILL10_259 <= 64'd0;
               Tsf1SPILL10_258 <= 64'd0;
               Tsin1_19_V_0 <= 32'd0;
               Tsin1_19_V_1 <= 32'd0;
               Tsco5_4_V_0 <= 32'd0;
               Tsco5_4_V_1 <= 32'd0;
               Tsin1_19_V_3 <= 32'd0;
               Tsin1_19_V_2 <= 64'd0;
               Tsi1_SPILL_256 <= 64'd0;
               Tsp5_SPILL_256 <= 64'd0;
               Tsi1_SPILL_257 <= 32'd0;
               Tsfl1_8_V_3 <= 32'd0;
               Tsfl1_8_V_4 <= 32'd0;
               Tsfl1_8_V_6 <= 64'd0;
               Tsfl1_8_V_7 <= 64'd0;
               fastspilldup28 <= 64'd0;
               fastspilldup30 <= 64'd0;
               Tsfl1_8_V_9 <= 64'd0;
               fastspilldup32 <= 64'd0;
               Tsf1_SPILL_260 <= 64'd0;
               Tsf1_SPILL_257 <= 64'd0;
               Tsfl1_8_V_8 <= 64'd0;
               Tsfl1_8_V_5 <= 32'd0;
               fastspilldup34 <= 64'd0;
               Tsf1_SPILL_256 <= 64'd0;
               fastspilldup36 <= 64'd0;
               Tsf1_SPILL_259 <= 64'd0;
               Tsf1_SPILL_258 <= 64'd0;
               Tsp4_SPILL_256 <= 64'd0;
               Tsp8_SPILL_256 <= 64'd0;
               Tspr11_2_V_2 <= 32'd0;
               Tspr11_2_V_3 <= 32'd0;
               Tspr11_2_V_4 <= 32'd0;
               Tspr11_2_V_0 <= 64'd0;
               Tspr11_2_V_1 <= 64'd0;
               Tsp11_SPILL_256 <= 64'd0;
               Tsf0SPILL12_256 <= 32'd0;
               Tsf0SPILL10_256 <= 32'd0;
               Tsp15_SPILL_256 <= 64'd0;
               Tsp18_SPILL_256 <= 64'd0;
               Tsno19_4_V_0 <= 32'd0;
               Tsfl0_9_V_3 <= 32'd0;
               Tsp22_SPILL_256 <= 64'd0;
               Tsco3_7_V_0 <= 32'd0;
               Tsco3_7_V_1 <= 32'd0;
               Tsco0_2_V_1 <= 32'd0;
               Tsno23_4_V_0 <= 32'd0;
               Tsfl0_9_V_4 <= 32'd0;
               Tsfl0_9_V_6 <= 64'd0;
               Tsfl0_9_V_7 <= 64'd0;
               Tsmu24_24_V_1 <= 32'd0;
               Tsmu24_24_V_0 <= 32'd0;
               Tsmu24_24_V_3 <= 32'd0;
               Tsmu24_24_V_2 <= 32'd0;
               Tsmu24_24_V_6 <= 64'd0;
               fastspilldup18 <= 64'd0;
               Tsm24_SPILL_264 <= 64'd0;
               Tsm24_SPILL_257 <= 64'd0;
               Tsmu24_24_V_5 <= 64'd0;
               Tsmu24_24_V_7 <= 64'd0;
               fastspilldup20 <= 64'd0;
               Tsm24_SPILL_263 <= 64'd0;
               Tsm24_SPILL_260 <= 64'd0;
               Tsmu24_24_V_4 <= 64'd0;
               Tsfl0_9_V_9 <= 64'd0;
               fastspilldup22 <= 64'd0;
               Tsf0_SPILL_260 <= 64'd0;
               Tsf0_SPILL_257 <= 64'd0;
               Tsfl0_9_V_8 <= 64'd0;
               Tsfl0_9_V_5 <= 32'd0;
               Tsro29_4_V_5 <= 32'd0;
               fastspilldup24 <= 64'd0;
               Tsr29_SPILL_260 <= 64'd0;
               Tsr29_SPILL_256 <= 64'd0;
               Tsf0_SPILL_256 <= 64'd0;
               Tsr29_SPILL_258 <= 64'd0;
               Tsr29_SPILL_257 <= 64'd0;
               Tsp13_SPILL_256 <= 64'd0;
               Tsro29_4_V_6 <= 32'd0;
               Tsro29_4_V_1 <= 64'd0;
               Tsro29_4_V_0 <= 32'd0;
               Tsr29_SPILL_259 <= 64'd0;
               Tsp27_SPILL_256 <= 64'd0;
               fastspilldup26 <= 64'd0;
               Tss18_SPILL_259 <= 64'd0;
               Tss18_SPILL_256 <= 64'd0;
               Tss18_SPILL_258 <= 64'd0;
               Tss18_SPILL_257 <= 64'd0;
               Tssh18_7_V_0 <= 64'd0;
               Tss18_SPILL_260 <= 64'd0;
               Tsf0_SPILL_259 <= 64'd0;
               Tsf0_SPILL_258 <= 64'd0;
               Tsm24_SPILL_262 <= 64'd0;
               Tsm24_SPILL_261 <= 64'd0;
               Tsm24_SPILL_259 <= 64'd0;
               Tsm24_SPILL_258 <= 64'd0;
               Tsco0_2_V_0 <= 64'd0;
               Tse0SPILL10_256 <= 32'd0;
               Tse0_SPILL_256 <= 32'd0;
               xpc10 <= 32'd0;
               end 
               else  begin 
              
              case (xpc10)
                  13'sd415/*415:xpc10*/: $display("dfsin: Testbench start");

                  13'sd515/*515:xpc10*/: $display("m_rad2=%H", Tdsi1_5_V_3);

                  13'sd520/*520:xpc10*/: $display("inc=%H", Tdsi1_5_V_2);

                  13'sd614/*614:xpc10*/: $display("nn=%H dd=%H", Tsf1_SPILL_256, Tsi1_SPILL_256);

                  13'sd872/*872:xpc10*/: $display(" diff=%H app=%H", Tdsi1_5_V_1, Tdsi1_5_V_0);

                  13'sd912/*912:xpc10*/: $display("Test: input=%H expected=%H output=%H ", A_64_US_CC_SCALbx12_ARB0[Tdbm0_3_V_1], A_64_US_CC_SCALbx10_ARA0
                  [Tdbm0_3_V_1], Tdbm0_3_V_2);

                  13'sd918/*918:xpc10*/: $display("   hamming error=%H", Tdbm0_3_V_2^A_64_US_CC_SCALbx10_ARA0[Tdbm0_3_V_1]);

                  13'sd932/*932:xpc10*/: $display("Result: %1d", Tdbm0_3_V_0);

                  13'sd938/*938:xpc10*/: $display("RESULT: PASS");

                  13'sd943/*943:xpc10*/: $display("dfsin: Testbench finished");
              endcase
              if ((13'sd948/*948:xpc10*/==xpc10)) $finish(32'sd0);
                  if ((13'sd951/*951:xpc10*/==xpc10)) $display("RESULT: FAIL");
                  if ((Tsco3_7_V_0<32'sh100_0000)) 
                  case (xpc10)
                      13'sd1727/*1727:xpc10*/:  xpc10 <= 13'sd1728/*1728:xpc10*/;

                      13'sd2544/*2544:xpc10*/:  xpc10 <= 13'sd2545/*2545:xpc10*/;

                      13'sd2606/*2606:xpc10*/:  xpc10 <= 13'sd2607/*2607:xpc10*/;

                      13'sd3382/*3382:xpc10*/:  xpc10 <= 13'sd3383/*3383:xpc10*/;

                      13'sd3444/*3444:xpc10*/:  xpc10 <= 13'sd3445/*3445:xpc10*/;

                      13'sd4004/*4004:xpc10*/:  xpc10 <= 13'sd4005/*4005:xpc10*/;

                      13'sd4066/*4066:xpc10*/:  xpc10 <= 13'sd4067/*4067:xpc10*/;

                      13'sd4573/*4573:xpc10*/:  xpc10 <= 13'sd4574/*4574:xpc10*/;

                      13'sd4635/*4635:xpc10*/:  xpc10 <= 13'sd4636/*4636:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd1727/*1727:xpc10*/:  xpc10 <= 13'sd1734/*1734:xpc10*/;

                      13'sd2544/*2544:xpc10*/:  xpc10 <= 13'sd2551/*2551:xpc10*/;

                      13'sd2606/*2606:xpc10*/:  xpc10 <= 13'sd2613/*2613:xpc10*/;

                      13'sd3382/*3382:xpc10*/:  xpc10 <= 13'sd3389/*3389:xpc10*/;

                      13'sd3444/*3444:xpc10*/:  xpc10 <= 13'sd3451/*3451:xpc10*/;

                      13'sd4004/*4004:xpc10*/:  xpc10 <= 13'sd4011/*4011:xpc10*/;

                      13'sd4066/*4066:xpc10*/:  xpc10 <= 13'sd4073/*4073:xpc10*/;

                      13'sd4573/*4573:xpc10*/:  xpc10 <= 13'sd4580/*4580:xpc10*/;

                      13'sd4635/*4635:xpc10*/:  xpc10 <= 13'sd4642/*4642:xpc10*/;
                  endcase
              if ((Tsco3_7_V_0<32'sh1_0000)) 
                  case (xpc10)
                      13'sd1718/*1718:xpc10*/:  xpc10 <= 13'sd1719/*1719:xpc10*/;

                      13'sd2535/*2535:xpc10*/:  xpc10 <= 13'sd2536/*2536:xpc10*/;

                      13'sd2597/*2597:xpc10*/:  xpc10 <= 13'sd2598/*2598:xpc10*/;

                      13'sd3373/*3373:xpc10*/:  xpc10 <= 13'sd3374/*3374:xpc10*/;

                      13'sd3435/*3435:xpc10*/:  xpc10 <= 13'sd3436/*3436:xpc10*/;

                      13'sd3995/*3995:xpc10*/:  xpc10 <= 13'sd3996/*3996:xpc10*/;

                      13'sd4057/*4057:xpc10*/:  xpc10 <= 13'sd4058/*4058:xpc10*/;

                      13'sd4564/*4564:xpc10*/:  xpc10 <= 13'sd4565/*4565:xpc10*/;

                      13'sd4626/*4626:xpc10*/:  xpc10 <= 13'sd4627/*4627:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd1718/*1718:xpc10*/:  xpc10 <= 13'sd1725/*1725:xpc10*/;

                      13'sd2535/*2535:xpc10*/:  xpc10 <= 13'sd2542/*2542:xpc10*/;

                      13'sd2597/*2597:xpc10*/:  xpc10 <= 13'sd2604/*2604:xpc10*/;

                      13'sd3373/*3373:xpc10*/:  xpc10 <= 13'sd3380/*3380:xpc10*/;

                      13'sd3435/*3435:xpc10*/:  xpc10 <= 13'sd3442/*3442:xpc10*/;

                      13'sd3995/*3995:xpc10*/:  xpc10 <= 13'sd4002/*4002:xpc10*/;

                      13'sd4057/*4057:xpc10*/:  xpc10 <= 13'sd4064/*4064:xpc10*/;

                      13'sd4564/*4564:xpc10*/:  xpc10 <= 13'sd4571/*4571:xpc10*/;

                      13'sd4626/*4626:xpc10*/:  xpc10 <= 13'sd4633/*4633:xpc10*/;
                  endcase
              if ((Tsco0_2_V_0<64'sh1_0000_0000)) 
                  case (xpc10)
                      13'sd1708/*1708:xpc10*/:  xpc10 <= 13'sd1709/*1709:xpc10*/;

                      13'sd2525/*2525:xpc10*/:  xpc10 <= 13'sd2526/*2526:xpc10*/;

                      13'sd2587/*2587:xpc10*/:  xpc10 <= 13'sd2588/*2588:xpc10*/;

                      13'sd3363/*3363:xpc10*/:  xpc10 <= 13'sd3364/*3364:xpc10*/;

                      13'sd3425/*3425:xpc10*/:  xpc10 <= 13'sd3426/*3426:xpc10*/;

                      13'sd3985/*3985:xpc10*/:  xpc10 <= 13'sd3986/*3986:xpc10*/;

                      13'sd4047/*4047:xpc10*/:  xpc10 <= 13'sd4048/*4048:xpc10*/;

                      13'sd4554/*4554:xpc10*/:  xpc10 <= 13'sd4555/*4555:xpc10*/;

                      13'sd4616/*4616:xpc10*/:  xpc10 <= 13'sd4617/*4617:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd1708/*1708:xpc10*/:  xpc10 <= 13'sd1909/*1909:xpc10*/;

                      13'sd2525/*2525:xpc10*/:  xpc10 <= 13'sd3105/*3105:xpc10*/;

                      13'sd2587/*2587:xpc10*/:  xpc10 <= 13'sd3101/*3101:xpc10*/;

                      13'sd3363/*3363:xpc10*/:  xpc10 <= 13'sd3727/*3727:xpc10*/;

                      13'sd3425/*3425:xpc10*/:  xpc10 <= 13'sd3723/*3723:xpc10*/;

                      13'sd3985/*3985:xpc10*/:  xpc10 <= 13'sd4349/*4349:xpc10*/;

                      13'sd4047/*4047:xpc10*/:  xpc10 <= 13'sd4345/*4345:xpc10*/;

                      13'sd4554/*4554:xpc10*/:  xpc10 <= 13'sd4918/*4918:xpc10*/;

                      13'sd4616/*4616:xpc10*/:  xpc10 <= 13'sd4914/*4914:xpc10*/;
                  endcase
              if (Tsfl0_9_V_2) 
                  case (xpc10)
                      13'sd4404/*4404:xpc10*/:  xpc10 <= 13'sd4405/*4405:xpc10*/;

                      13'sd4512/*4512:xpc10*/:  xpc10 <= 13'sd4513/*4513:xpc10*/;

                      13'sd4536/*4536:xpc10*/:  xpc10 <= 13'sd4537/*4537:xpc10*/;

                      13'sd4598/*4598:xpc10*/:  xpc10 <= 13'sd4599/*4599:xpc10*/;

                      13'sd4751/*4751:xpc10*/:  xpc10 <= 13'sd4752/*4752:xpc10*/;

                      13'sd4840/*4840:xpc10*/:  xpc10 <= 13'sd4841/*4841:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd4404/*4404:xpc10*/:  xpc10 <= 13'sd4414/*4414:xpc10*/;

                      13'sd4512/*4512:xpc10*/:  xpc10 <= 13'sd4522/*4522:xpc10*/;

                      13'sd4536/*4536:xpc10*/:  xpc10 <= 13'sd4546/*4546:xpc10*/;

                      13'sd4598/*4598:xpc10*/:  xpc10 <= 13'sd4608/*4608:xpc10*/;

                      13'sd4751/*4751:xpc10*/:  xpc10 <= 13'sd4782/*4782:xpc10*/;

                      13'sd4840/*4840:xpc10*/:  xpc10 <= 13'sd4850/*4850:xpc10*/;
                  endcase
              if (Tsfl1_8_V_2) 
                  case (xpc10)
                      13'sd3835/*3835:xpc10*/:  xpc10 <= 13'sd3836/*3836:xpc10*/;

                      13'sd3943/*3943:xpc10*/:  xpc10 <= 13'sd3944/*3944:xpc10*/;

                      13'sd3967/*3967:xpc10*/:  xpc10 <= 13'sd3968/*3968:xpc10*/;

                      13'sd4029/*4029:xpc10*/:  xpc10 <= 13'sd4030/*4030:xpc10*/;

                      13'sd4182/*4182:xpc10*/:  xpc10 <= 13'sd4183/*4183:xpc10*/;

                      13'sd4271/*4271:xpc10*/:  xpc10 <= 13'sd4272/*4272:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd3835/*3835:xpc10*/:  xpc10 <= 13'sd3845/*3845:xpc10*/;

                      13'sd3943/*3943:xpc10*/:  xpc10 <= 13'sd3953/*3953:xpc10*/;

                      13'sd3967/*3967:xpc10*/:  xpc10 <= 13'sd3977/*3977:xpc10*/;

                      13'sd4029/*4029:xpc10*/:  xpc10 <= 13'sd4039/*4039:xpc10*/;

                      13'sd4182/*4182:xpc10*/:  xpc10 <= 13'sd4213/*4213:xpc10*/;

                      13'sd4271/*4271:xpc10*/:  xpc10 <= 13'sd4281/*4281:xpc10*/;
                  endcase
              if ((Tsro29_4_V_1==32'sd0/*0:Tsro29.4_V_1*/)) 
                  case (xpc10)
                      13'sd3641/*3641:xpc10*/:  xpc10 <= 13'sd3642/*3642:xpc10*/;

                      13'sd3690/*3690:xpc10*/:  xpc10 <= 13'sd3700/*3700:xpc10*/;

                      13'sd4263/*4263:xpc10*/:  xpc10 <= 13'sd4264/*4264:xpc10*/;

                      13'sd4312/*4312:xpc10*/:  xpc10 <= 13'sd4322/*4322:xpc10*/;

                      13'sd4832/*4832:xpc10*/:  xpc10 <= 13'sd4833/*4833:xpc10*/;

                      13'sd4881/*4881:xpc10*/:  xpc10 <= 13'sd4891/*4891:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd3641/*3641:xpc10*/:  xpc10 <= 13'sd3647/*3647:xpc10*/;

                      13'sd3690/*3690:xpc10*/:  xpc10 <= 13'sd3691/*3691:xpc10*/;

                      13'sd4263/*4263:xpc10*/:  xpc10 <= 13'sd4269/*4269:xpc10*/;

                      13'sd4312/*4312:xpc10*/:  xpc10 <= 13'sd4313/*4313:xpc10*/;

                      13'sd4832/*4832:xpc10*/:  xpc10 <= 13'sd4838/*4838:xpc10*/;

                      13'sd4881/*4881:xpc10*/:  xpc10 <= 13'sd4882/*4882:xpc10*/;
                  endcase
              if (!(!Tsro29_4_V_6)) 
                  case (xpc10)
                      13'sd3616/*3616:xpc10*/:  xpc10 <= 13'sd3617/*3617:xpc10*/;

                      13'sd3624/*3624:xpc10*/:  xpc10 <= 13'sd3625/*3625:xpc10*/;

                      13'sd4238/*4238:xpc10*/:  xpc10 <= 13'sd4239/*4239:xpc10*/;

                      13'sd4246/*4246:xpc10*/:  xpc10 <= 13'sd4247/*4247:xpc10*/;

                      13'sd4807/*4807:xpc10*/:  xpc10 <= 13'sd4808/*4808:xpc10*/;

                      13'sd4815/*4815:xpc10*/:  xpc10 <= 13'sd4816/*4816:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd3616/*3616:xpc10*/:  xpc10 <= 13'sd3622/*3622:xpc10*/;

                      13'sd3624/*3624:xpc10*/:  xpc10 <= 13'sd3630/*3630:xpc10*/;

                      13'sd4238/*4238:xpc10*/:  xpc10 <= 13'sd4244/*4244:xpc10*/;

                      13'sd4246/*4246:xpc10*/:  xpc10 <= 13'sd4252/*4252:xpc10*/;

                      13'sd4807/*4807:xpc10*/:  xpc10 <= 13'sd4813/*4813:xpc10*/;

                      13'sd4815/*4815:xpc10*/:  xpc10 <= 13'sd4821/*4821:xpc10*/;
                  endcase
              if ((Tsmu24_24_V_5<Tsmu24_24_V_6)) 
                  case (xpc10)
                      13'sd3473/*3473:xpc10*/:  xpc10 <= 13'sd3474/*3474:xpc10*/;

                      13'sd3485/*3485:xpc10*/:  xpc10 <= 13'sd3486/*3486:xpc10*/;

                      13'sd4095/*4095:xpc10*/:  xpc10 <= 13'sd4096/*4096:xpc10*/;

                      13'sd4107/*4107:xpc10*/:  xpc10 <= 13'sd4108/*4108:xpc10*/;

                      13'sd4664/*4664:xpc10*/:  xpc10 <= 13'sd4665/*4665:xpc10*/;

                      13'sd4676/*4676:xpc10*/:  xpc10 <= 13'sd4677/*4677:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd3473/*3473:xpc10*/:  xpc10 <= 13'sd3719/*3719:xpc10*/;

                      13'sd3485/*3485:xpc10*/:  xpc10 <= 13'sd3714/*3714:xpc10*/;

                      13'sd4095/*4095:xpc10*/:  xpc10 <= 13'sd4341/*4341:xpc10*/;

                      13'sd4107/*4107:xpc10*/:  xpc10 <= 13'sd4336/*4336:xpc10*/;

                      13'sd4664/*4664:xpc10*/:  xpc10 <= 13'sd4910/*4910:xpc10*/;

                      13'sd4676/*4676:xpc10*/:  xpc10 <= 13'sd4905/*4905:xpc10*/;
                  endcase
              if (Tsfl1_24_V_2) 
                  case (xpc10)
                      13'sd3213/*3213:xpc10*/:  xpc10 <= 13'sd3214/*3214:xpc10*/;

                      13'sd3321/*3321:xpc10*/:  xpc10 <= 13'sd3322/*3322:xpc10*/;

                      13'sd3345/*3345:xpc10*/:  xpc10 <= 13'sd3346/*3346:xpc10*/;

                      13'sd3407/*3407:xpc10*/:  xpc10 <= 13'sd3408/*3408:xpc10*/;

                      13'sd3560/*3560:xpc10*/:  xpc10 <= 13'sd3561/*3561:xpc10*/;

                      13'sd3649/*3649:xpc10*/:  xpc10 <= 13'sd3650/*3650:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd3213/*3213:xpc10*/:  xpc10 <= 13'sd3223/*3223:xpc10*/;

                      13'sd3321/*3321:xpc10*/:  xpc10 <= 13'sd3331/*3331:xpc10*/;

                      13'sd3345/*3345:xpc10*/:  xpc10 <= 13'sd3355/*3355:xpc10*/;

                      13'sd3407/*3407:xpc10*/:  xpc10 <= 13'sd3417/*3417:xpc10*/;

                      13'sd3560/*3560:xpc10*/:  xpc10 <= 13'sd3591/*3591:xpc10*/;

                      13'sd3649/*3649:xpc10*/:  xpc10 <= 13'sd3659/*3659:xpc10*/;
                  endcase
              if (Tsfl1_35_V_2) 
                  case (xpc10)
                      13'sd2374/*2374:xpc10*/:  xpc10 <= 13'sd2375/*2375:xpc10*/;

                      13'sd2469/*2469:xpc10*/:  xpc10 <= 13'sd2470/*2470:xpc10*/;

                      13'sd2507/*2507:xpc10*/:  xpc10 <= 13'sd2508/*2508:xpc10*/;

                      13'sd2569/*2569:xpc10*/:  xpc10 <= 13'sd2570/*2570:xpc10*/;

                      13'sd2759/*2759:xpc10*/:  xpc10 <= 13'sd2760/*2760:xpc10*/;

                      13'sd2848/*2848:xpc10*/:  xpc10 <= 13'sd2849/*2849:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd2374/*2374:xpc10*/:  xpc10 <= 13'sd2384/*2384:xpc10*/;

                      13'sd2469/*2469:xpc10*/:  xpc10 <= 13'sd2479/*2479:xpc10*/;

                      13'sd2507/*2507:xpc10*/:  xpc10 <= 13'sd2517/*2517:xpc10*/;

                      13'sd2569/*2569:xpc10*/:  xpc10 <= 13'sd2579/*2579:xpc10*/;

                      13'sd2759/*2759:xpc10*/:  xpc10 <= 13'sd2790/*2790:xpc10*/;

                      13'sd2848/*2848:xpc10*/:  xpc10 <= 13'sd2858/*2858:xpc10*/;
                  endcase
              if (Tsfl1_39_V_0) 
                  case (xpc10)
                      13'sd1109/*1109:xpc10*/:  xpc10 <= 13'sd1110/*1110:xpc10*/;

                      13'sd1198/*1198:xpc10*/:  xpc10 <= 13'sd1199/*1199:xpc10*/;

                      13'sd1383/*1383:xpc10*/:  xpc10 <= 13'sd1384/*1384:xpc10*/;

                      13'sd1556/*1556:xpc10*/:  xpc10 <= 13'sd1557/*1557:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd1109/*1109:xpc10*/:  xpc10 <= 13'sd1140/*1140:xpc10*/;

                      13'sd1198/*1198:xpc10*/:  xpc10 <= 13'sd1208/*1208:xpc10*/;

                      13'sd1383/*1383:xpc10*/:  xpc10 <= 13'sd1393/*1393:xpc10*/;

                      13'sd1556/*1556:xpc10*/:  xpc10 <= 13'sd1566/*1566:xpc10*/;
                  endcase
              if ((Tsfl1_24_V_7==32'sd0/*0:Tsfl1.24_V_7*/)) 
                  case (xpc10)
                      13'sd653/*653:xpc10*/:  xpc10 <= 13'sd3198/*3198:xpc10*/;

                      13'sd3204/*3204:xpc10*/:  xpc10 <= 13'sd3205/*3205:xpc10*/;

                      13'sd3233/*3233:xpc10*/:  xpc10 <= 13'sd3306/*3306:xpc10*/;

                      13'sd3403/*3403:xpc10*/:  xpc10 <= 13'sd3404/*3404:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd653/*653:xpc10*/:  xpc10 <= 13'sd654/*654:xpc10*/;

                      13'sd3204/*3204:xpc10*/:  xpc10 <= 13'sd3211/*3211:xpc10*/;

                      13'sd3233/*3233:xpc10*/:  xpc10 <= 13'sd3234/*3234:xpc10*/;

                      13'sd3403/*3403:xpc10*/:  xpc10 <= 13'sd3421/*3421:xpc10*/;
                  endcase
              if ((Tsfl1_8_V_7==32'sd0/*0:Tsfl1.8_V_7*/)) 
                  case (xpc10)
                      13'sd559/*559:xpc10*/:  xpc10 <= 13'sd3820/*3820:xpc10*/;

                      13'sd3826/*3826:xpc10*/:  xpc10 <= 13'sd3827/*3827:xpc10*/;

                      13'sd3855/*3855:xpc10*/:  xpc10 <= 13'sd3928/*3928:xpc10*/;

                      13'sd4025/*4025:xpc10*/:  xpc10 <= 13'sd4026/*4026:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd559/*559:xpc10*/:  xpc10 <= 13'sd560/*560:xpc10*/;

                      13'sd3826/*3826:xpc10*/:  xpc10 <= 13'sd3833/*3833:xpc10*/;

                      13'sd3855/*3855:xpc10*/:  xpc10 <= 13'sd3856/*3856:xpc10*/;

                      13'sd4025/*4025:xpc10*/:  xpc10 <= 13'sd4043/*4043:xpc10*/;
                  endcase
              if ((Tsfl0_9_V_7==32'sd0/*0:Tsfl0.9_V_7*/)) 
                  case (xpc10)
                      13'sd466/*466:xpc10*/:  xpc10 <= 13'sd4389/*4389:xpc10*/;

                      13'sd4395/*4395:xpc10*/:  xpc10 <= 13'sd4396/*4396:xpc10*/;

                      13'sd4424/*4424:xpc10*/:  xpc10 <= 13'sd4497/*4497:xpc10*/;

                      13'sd4594/*4594:xpc10*/:  xpc10 <= 13'sd4595/*4595:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd466/*466:xpc10*/:  xpc10 <= 13'sd467/*467:xpc10*/;

                      13'sd4395/*4395:xpc10*/:  xpc10 <= 13'sd4402/*4402:xpc10*/;

                      13'sd4424/*4424:xpc10*/:  xpc10 <= 13'sd4425/*4425:xpc10*/;

                      13'sd4594/*4594:xpc10*/:  xpc10 <= 13'sd4612/*4612:xpc10*/;
                  endcase
              if ((32'sd0/*0:USA34*/==(Tsro29_4_V_1<<(32'sd63&rtl_signed_bitextract0(Tsro29_4_V_0))))) 
                  case (xpc10)
                      13'sd3672/*3672:xpc10*/:  xpc10 <= 13'sd3683/*3683:xpc10*/;

                      13'sd4294/*4294:xpc10*/:  xpc10 <= 13'sd4305/*4305:xpc10*/;

                      13'sd4863/*4863:xpc10*/:  xpc10 <= 13'sd4874/*4874:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd3672/*3672:xpc10*/:  xpc10 <= 13'sd3673/*3673:xpc10*/;

                      13'sd4294/*4294:xpc10*/:  xpc10 <= 13'sd4295/*4295:xpc10*/;

                      13'sd4863/*4863:xpc10*/:  xpc10 <= 13'sd4864/*4864:xpc10*/;
                  endcase
              if ((rtl_signed_bitextract0((0-Tsro29_4_V_0))<32'sd64)) 
                  case (xpc10)
                      13'sd3665/*3665:xpc10*/:  xpc10 <= 13'sd3666/*3666:xpc10*/;

                      13'sd4287/*4287:xpc10*/:  xpc10 <= 13'sd4288/*4288:xpc10*/;

                      13'sd4856/*4856:xpc10*/:  xpc10 <= 13'sd4857/*4857:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd3665/*3665:xpc10*/:  xpc10 <= 13'sd3688/*3688:xpc10*/;

                      13'sd4287/*4287:xpc10*/:  xpc10 <= 13'sd4310/*4310:xpc10*/;

                      13'sd4856/*4856:xpc10*/:  xpc10 <= 13'sd4879/*4879:xpc10*/;
                  endcase
              if (32'sd1&(32'sd0/*0:USA36*/==(32'sd512^Tsro29_4_V_6))) 
                  case (xpc10)
                      13'sd3633/*3633:xpc10*/:  xpc10 <= 13'sd3634/*3634:xpc10*/;

                      13'sd4255/*4255:xpc10*/:  xpc10 <= 13'sd4256/*4256:xpc10*/;

                      13'sd4824/*4824:xpc10*/:  xpc10 <= 13'sd4825/*4825:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd3633/*3633:xpc10*/:  xpc10 <= 13'sd3639/*3639:xpc10*/;

                      13'sd4255/*4255:xpc10*/:  xpc10 <= 13'sd4261/*4261:xpc10*/;

                      13'sd4824/*4824:xpc10*/:  xpc10 <= 13'sd4830/*4830:xpc10*/;
                  endcase
              if (!(!rtl_signed_bitextract0((0-Tsro29_4_V_0)))) 
                  case (xpc10)
                      13'sd3602/*3602:xpc10*/:  xpc10 <= 13'sd3663/*3663:xpc10*/;

                      13'sd4224/*4224:xpc10*/:  xpc10 <= 13'sd4285/*4285:xpc10*/;

                      13'sd4793/*4793:xpc10*/:  xpc10 <= 13'sd4854/*4854:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd3602/*3602:xpc10*/:  xpc10 <= 13'sd3603/*3603:xpc10*/;

                      13'sd4224/*4224:xpc10*/:  xpc10 <= 13'sd4225/*4225:xpc10*/;

                      13'sd4793/*4793:xpc10*/:  xpc10 <= 13'sd4794/*4794:xpc10*/;
                  endcase
              if ((Tsro29_4_V_0<32'sd0)) 
                  case (xpc10)
                      13'sd3597/*3597:xpc10*/:  xpc10 <= 13'sd3598/*3598:xpc10*/;

                      13'sd4219/*4219:xpc10*/:  xpc10 <= 13'sd4220/*4220:xpc10*/;

                      13'sd4788/*4788:xpc10*/:  xpc10 <= 13'sd4789/*4789:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd3597/*3597:xpc10*/:  xpc10 <= 13'sd3622/*3622:xpc10*/;

                      13'sd4219/*4219:xpc10*/:  xpc10 <= 13'sd4244/*4244:xpc10*/;

                      13'sd4788/*4788:xpc10*/:  xpc10 <= 13'sd4813/*4813:xpc10*/;
                  endcase
              if (!(!Tsro29_4_V_5)) 
                  case (xpc10)
                      13'sd3571/*3571:xpc10*/:  xpc10 <= 13'sd3586/*3586:xpc10*/;

                      13'sd4193/*4193:xpc10*/:  xpc10 <= 13'sd4208/*4208:xpc10*/;

                      13'sd4762/*4762:xpc10*/:  xpc10 <= 13'sd4777/*4777:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd3571/*3571:xpc10*/:  xpc10 <= 13'sd3572/*3572:xpc10*/;

                      13'sd4193/*4193:xpc10*/:  xpc10 <= 13'sd4194/*4194:xpc10*/;

                      13'sd4762/*4762:xpc10*/:  xpc10 <= 13'sd4763/*4763:xpc10*/;
                  endcase
              if ((Tsro29_4_V_1+rtl_sign_extend1(Tsro29_4_V_5)<64'sh0)) 
                  case (xpc10)
                      13'sd3555/*3555:xpc10*/:  xpc10 <= 13'sd3556/*3556:xpc10*/;

                      13'sd4177/*4177:xpc10*/:  xpc10 <= 13'sd4178/*4178:xpc10*/;

                      13'sd4746/*4746:xpc10*/:  xpc10 <= 13'sd4747/*4747:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd3555/*3555:xpc10*/:  xpc10 <= 13'sd3595/*3595:xpc10*/;

                      13'sd4177/*4177:xpc10*/:  xpc10 <= 13'sd4217/*4217:xpc10*/;

                      13'sd4746/*4746:xpc10*/:  xpc10 <= 13'sd4786/*4786:xpc10*/;
                  endcase
              if ((Tsro29_4_V_0==32'sd2045/*2045:Tsro29.4_V_0*/)) 
                  case (xpc10)
                      13'sd3551/*3551:xpc10*/:  xpc10 <= 13'sd3552/*3552:xpc10*/;

                      13'sd4173/*4173:xpc10*/:  xpc10 <= 13'sd4174/*4174:xpc10*/;

                      13'sd4742/*4742:xpc10*/:  xpc10 <= 13'sd4743/*4743:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd3551/*3551:xpc10*/:  xpc10 <= 13'sd3595/*3595:xpc10*/;

                      13'sd4173/*4173:xpc10*/:  xpc10 <= 13'sd4217/*4217:xpc10*/;

                      13'sd4742/*4742:xpc10*/:  xpc10 <= 13'sd4786/*4786:xpc10*/;
                  endcase
              if ((32'sd2045<Tsro29_4_V_0)) 
                  case (xpc10)
                      13'sd3547/*3547:xpc10*/:  xpc10 <= 13'sd3557/*3557:xpc10*/;

                      13'sd4169/*4169:xpc10*/:  xpc10 <= 13'sd4179/*4179:xpc10*/;

                      13'sd4738/*4738:xpc10*/:  xpc10 <= 13'sd4748/*4748:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd3547/*3547:xpc10*/:  xpc10 <= 13'sd3548/*3548:xpc10*/;

                      13'sd4169/*4169:xpc10*/:  xpc10 <= 13'sd4170/*4170:xpc10*/;

                      13'sd4738/*4738:xpc10*/:  xpc10 <= 13'sd4739/*4739:xpc10*/;
                  endcase
              if ((Tsro29_4_V_0<32'sd2045)) 
                  case (xpc10)
                      13'sd3543/*3543:xpc10*/:  xpc10 <= 13'sd3622/*3622:xpc10*/;

                      13'sd4165/*4165:xpc10*/:  xpc10 <= 13'sd4244/*4244:xpc10*/;

                      13'sd4734/*4734:xpc10*/:  xpc10 <= 13'sd4813/*4813:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd3543/*3543:xpc10*/:  xpc10 <= 13'sd3544/*3544:xpc10*/;

                      13'sd4165/*4165:xpc10*/:  xpc10 <= 13'sd4166/*4166:xpc10*/;

                      13'sd4734/*4734:xpc10*/:  xpc10 <= 13'sd4735/*4735:xpc10*/;
                  endcase
              if ((Tsmu24_24_V_7<Tsmu24_24_V_5)) 
                  case (xpc10)
                      13'sd3500/*3500:xpc10*/:  xpc10 <= 13'sd3501/*3501:xpc10*/;

                      13'sd4122/*4122:xpc10*/:  xpc10 <= 13'sd4123/*4123:xpc10*/;

                      13'sd4691/*4691:xpc10*/:  xpc10 <= 13'sd4692/*4692:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd3500/*3500:xpc10*/:  xpc10 <= 13'sd3709/*3709:xpc10*/;

                      13'sd4122/*4122:xpc10*/:  xpc10 <= 13'sd4331/*4331:xpc10*/;

                      13'sd4691/*4691:xpc10*/:  xpc10 <= 13'sd4900/*4900:xpc10*/;
                  endcase
              if (Tspr11_2_V_3) 
                  case (xpc10)
                      13'sd3288/*3288:xpc10*/:  xpc10 <= 13'sd3289/*3289:xpc10*/;

                      13'sd3910/*3910:xpc10*/:  xpc10 <= 13'sd3911/*3911:xpc10*/;

                      13'sd4479/*4479:xpc10*/:  xpc10 <= 13'sd4480/*4480:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd3288/*3288:xpc10*/:  xpc10 <= 13'sd3294/*3294:xpc10*/;

                      13'sd3910/*3910:xpc10*/:  xpc10 <= 13'sd3916/*3916:xpc10*/;

                      13'sd4479/*4479:xpc10*/:  xpc10 <= 13'sd4485/*4485:xpc10*/;
                  endcase
              if (Tspr11_2_V_2) 
                  case (xpc10)
                      13'sd3280/*3280:xpc10*/:  xpc10 <= 13'sd3281/*3281:xpc10*/;

                      13'sd3902/*3902:xpc10*/:  xpc10 <= 13'sd3903/*3903:xpc10*/;

                      13'sd4471/*4471:xpc10*/:  xpc10 <= 13'sd4472/*4472:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd3280/*3280:xpc10*/:  xpc10 <= 13'sd3286/*3286:xpc10*/;

                      13'sd3902/*3902:xpc10*/:  xpc10 <= 13'sd3908/*3908:xpc10*/;

                      13'sd4471/*4471:xpc10*/:  xpc10 <= 13'sd4477/*4477:xpc10*/;
                  endcase
              if (Tspr11_2_V_4) 
                  case (xpc10)
                      13'sd3268/*3268:xpc10*/:  xpc10 <= 13'sd3269/*3269:xpc10*/;

                      13'sd3890/*3890:xpc10*/:  xpc10 <= 13'sd3891/*3891:xpc10*/;

                      13'sd4459/*4459:xpc10*/:  xpc10 <= 13'sd4460/*4460:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd3268/*3268:xpc10*/:  xpc10 <= 13'sd3278/*3278:xpc10*/;

                      13'sd3890/*3890:xpc10*/:  xpc10 <= 13'sd3900/*3900:xpc10*/;

                      13'sd4459/*4459:xpc10*/:  xpc10 <= 13'sd4469/*4469:xpc10*/;
                  endcase
              if ((32'sd4094/*4094:USA28*/==(64'shfff&(Tspr11_2_V_1>>32'sd51)))) 
                  case (xpc10)
                      13'sd3249/*3249:xpc10*/:  xpc10 <= 13'sd3250/*3250:xpc10*/;

                      13'sd3871/*3871:xpc10*/:  xpc10 <= 13'sd3872/*3872:xpc10*/;

                      13'sd4440/*4440:xpc10*/:  xpc10 <= 13'sd4441/*4441:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd3249/*3249:xpc10*/:  xpc10 <= 13'sd3298/*3298:xpc10*/;

                      13'sd3871/*3871:xpc10*/:  xpc10 <= 13'sd3920/*3920:xpc10*/;

                      13'sd4440/*4440:xpc10*/:  xpc10 <= 13'sd4489/*4489:xpc10*/;
                  endcase
              if ((32'sd4094/*4094:USA22*/==(64'shfff&(Tspr11_2_V_0>>32'sd51)))) 
                  case (xpc10)
                      13'sd3239/*3239:xpc10*/:  xpc10 <= 13'sd3240/*3240:xpc10*/;

                      13'sd3861/*3861:xpc10*/:  xpc10 <= 13'sd3862/*3862:xpc10*/;

                      13'sd4430/*4430:xpc10*/:  xpc10 <= 13'sd4431/*4431:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd3239/*3239:xpc10*/:  xpc10 <= 13'sd3302/*3302:xpc10*/;

                      13'sd3861/*3861:xpc10*/:  xpc10 <= 13'sd3924/*3924:xpc10*/;

                      13'sd4430/*4430:xpc10*/:  xpc10 <= 13'sd4493/*4493:xpc10*/;
                  endcase
              if (Tspr4_3_V_3) 
                  case (xpc10)
                      13'sd3180/*3180:xpc10*/:  xpc10 <= 13'sd3181/*3181:xpc10*/;

                      13'sd3802/*3802:xpc10*/:  xpc10 <= 13'sd3803/*3803:xpc10*/;

                      13'sd4371/*4371:xpc10*/:  xpc10 <= 13'sd4372/*4372:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd3180/*3180:xpc10*/:  xpc10 <= 13'sd3186/*3186:xpc10*/;

                      13'sd3802/*3802:xpc10*/:  xpc10 <= 13'sd3808/*3808:xpc10*/;

                      13'sd4371/*4371:xpc10*/:  xpc10 <= 13'sd4377/*4377:xpc10*/;
                  endcase
              if (Tspr4_3_V_2) 
                  case (xpc10)
                      13'sd3172/*3172:xpc10*/:  xpc10 <= 13'sd3173/*3173:xpc10*/;

                      13'sd3794/*3794:xpc10*/:  xpc10 <= 13'sd3795/*3795:xpc10*/;

                      13'sd4363/*4363:xpc10*/:  xpc10 <= 13'sd4364/*4364:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd3172/*3172:xpc10*/:  xpc10 <= 13'sd3178/*3178:xpc10*/;

                      13'sd3794/*3794:xpc10*/:  xpc10 <= 13'sd3800/*3800:xpc10*/;

                      13'sd4363/*4363:xpc10*/:  xpc10 <= 13'sd4369/*4369:xpc10*/;
                  endcase
              if ((Tsfl1_35_V_7==32'sd0/*0:Tsfl1.35_V_7*/)) 
                  case (xpc10)
                      13'sd2294/*2294:xpc10*/:  xpc10 <= 13'sd2367/*2367:xpc10*/;

                      13'sd2394/*2394:xpc10*/:  xpc10 <= 13'sd2467/*2467:xpc10*/;

                      13'sd2489/*2489:xpc10*/:  xpc10 <= 13'sd2490/*2490:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd2294/*2294:xpc10*/:  xpc10 <= 13'sd2295/*2295:xpc10*/;

                      13'sd2394/*2394:xpc10*/:  xpc10 <= 13'sd2395/*2395:xpc10*/;

                      13'sd2489/*2489:xpc10*/:  xpc10 <= 13'sd2521/*2521:xpc10*/;
                  endcase
              if ((Tssu2_4_V_5==32'sd0/*0:Tssu2.4_V_5*/)) 
                  case (xpc10)
                      13'sd1940/*1940:xpc10*/:  xpc10 <= 13'sd1950/*1950:xpc10*/;

                      13'sd1971/*1971:xpc10*/:  xpc10 <= 13'sd2044/*2044:xpc10*/;

                      13'sd2142/*2142:xpc10*/:  xpc10 <= 13'sd2215/*2215:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd1940/*1940:xpc10*/:  xpc10 <= 13'sd1941/*1941:xpc10*/;

                      13'sd1971/*1971:xpc10*/:  xpc10 <= 13'sd1972/*1972:xpc10*/;

                      13'sd2142/*2142:xpc10*/:  xpc10 <= 13'sd2143/*2143:xpc10*/;
                  endcase
              if ((Tssu2_4_V_4==32'sd0/*0:Tssu2.4_V_4*/)) 
                  case (xpc10)
                      13'sd1596/*1596:xpc10*/:  xpc10 <= 13'sd1673/*1673:xpc10*/;

                      13'sd2114/*2114:xpc10*/:  xpc10 <= 13'sd2124/*2124:xpc10*/;

                      13'sd2138/*2138:xpc10*/:  xpc10 <= 13'sd2139/*2139:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd1596/*1596:xpc10*/:  xpc10 <= 13'sd1597/*1597:xpc10*/;

                      13'sd2114/*2114:xpc10*/:  xpc10 <= 13'sd2115/*2115:xpc10*/;

                      13'sd2138/*2138:xpc10*/:  xpc10 <= 13'sd2144/*2144:xpc10*/;
                  endcase
              if ((Tsad1_3_V_4==32'sd0/*0:Tsad1.3_V_4*/)) 
                  case (xpc10)
                      13'sd1280/*1280:xpc10*/:  xpc10 <= 13'sd1290/*1290:xpc10*/;

                      13'sd1308/*1308:xpc10*/:  xpc10 <= 13'sd1381/*1381:xpc10*/;

                      13'sd1473/*1473:xpc10*/:  xpc10 <= 13'sd1546/*1546:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd1280/*1280:xpc10*/:  xpc10 <= 13'sd1281/*1281:xpc10*/;

                      13'sd1308/*1308:xpc10*/:  xpc10 <= 13'sd1309/*1309:xpc10*/;

                      13'sd1473/*1473:xpc10*/:  xpc10 <= 13'sd1474/*1474:xpc10*/;
                  endcase
              if ((Tsad1_3_V_3==32'sd0/*0:Tsad1.3_V_3*/)) 
                  case (xpc10)
                      13'sd820/*820:xpc10*/:  xpc10 <= 13'sd1044/*1044:xpc10*/;

                      13'sd1445/*1445:xpc10*/:  xpc10 <= 13'sd1455/*1455:xpc10*/;

                      13'sd1469/*1469:xpc10*/:  xpc10 <= 13'sd1470/*1470:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd820/*820:xpc10*/:  xpc10 <= 13'sd821/*821:xpc10*/;

                      13'sd1445/*1445:xpc10*/:  xpc10 <= 13'sd1446/*1446:xpc10*/;

                      13'sd1469/*1469:xpc10*/:  xpc10 <= 13'sd1475/*1475:xpc10*/;
                  endcase
              if ((Tsfl1_35_V_6==32'sd0/*0:Tsfl1.35_V_6*/)) 
                  case (xpc10)
                      13'sd735/*735:xpc10*/:  xpc10 <= 13'sd2288/*2288:xpc10*/;

                      13'sd2497/*2497:xpc10*/:  xpc10 <= 13'sd2498/*2498:xpc10*/;

                      13'sd2565/*2565:xpc10*/:  xpc10 <= 13'sd2566/*2566:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd735/*735:xpc10*/:  xpc10 <= 13'sd736/*736:xpc10*/;

                      13'sd2497/*2497:xpc10*/:  xpc10 <= 13'sd2504/*2504:xpc10*/;

                      13'sd2565/*2565:xpc10*/:  xpc10 <= 13'sd2583/*2583:xpc10*/;
                  endcase
              if ((Tsfl1_24_V_6==32'sd0/*0:Tsfl1.24_V_6*/)) 
                  case (xpc10)
                      13'sd645/*645:xpc10*/:  xpc10 <= 13'sd646/*646:xpc10*/;

                      13'sd3312/*3312:xpc10*/:  xpc10 <= 13'sd3313/*3313:xpc10*/;

                      13'sd3341/*3341:xpc10*/:  xpc10 <= 13'sd3342/*3342:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd645/*645:xpc10*/:  xpc10 <= 13'sd655/*655:xpc10*/;

                      13'sd3312/*3312:xpc10*/:  xpc10 <= 13'sd3319/*3319:xpc10*/;

                      13'sd3341/*3341:xpc10*/:  xpc10 <= 13'sd3359/*3359:xpc10*/;
                  endcase
              if ((Tsfl1_8_V_6==32'sd0/*0:Tsfl1.8_V_6*/)) 
                  case (xpc10)
                      13'sd551/*551:xpc10*/:  xpc10 <= 13'sd552/*552:xpc10*/;

                      13'sd3934/*3934:xpc10*/:  xpc10 <= 13'sd3935/*3935:xpc10*/;

                      13'sd3963/*3963:xpc10*/:  xpc10 <= 13'sd3964/*3964:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd551/*551:xpc10*/:  xpc10 <= 13'sd561/*561:xpc10*/;

                      13'sd3934/*3934:xpc10*/:  xpc10 <= 13'sd3941/*3941:xpc10*/;

                      13'sd3963/*3963:xpc10*/:  xpc10 <= 13'sd3981/*3981:xpc10*/;
                  endcase
              if ((64'sh0<(Tdsi1_5_V_1>>32'sd63))) 
                  case (xpc10)
                      13'sd526/*526:xpc10*/:  xpc10 <= 13'sd527/*527:xpc10*/;

                      13'sd620/*620:xpc10*/:  xpc10 <= 13'sd621/*621:xpc10*/;

                      13'sd792/*792:xpc10*/:  xpc10 <= 13'sd793/*793:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd526/*526:xpc10*/:  xpc10 <= 13'sd4357/*4357:xpc10*/;

                      13'sd620/*620:xpc10*/:  xpc10 <= 13'sd3735/*3735:xpc10*/;

                      13'sd792/*792:xpc10*/:  xpc10 <= 13'sd2252/*2252:xpc10*/;
                  endcase
              if (Tspr4_3_V_4) 
                  case (xpc10)
                      13'sd501/*501:xpc10*/:  xpc10 <= 13'sd502/*502:xpc10*/;

                      13'sd594/*594:xpc10*/:  xpc10 <= 13'sd595/*595:xpc10*/;

                      13'sd688/*688:xpc10*/:  xpc10 <= 13'sd689/*689:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd501/*501:xpc10*/:  xpc10 <= 13'sd4361/*4361:xpc10*/;

                      13'sd594/*594:xpc10*/:  xpc10 <= 13'sd3792/*3792:xpc10*/;

                      13'sd688/*688:xpc10*/:  xpc10 <= 13'sd3170/*3170:xpc10*/;
                  endcase
              if ((32'sd4094/*4094:USA16*/==(64'shfff&(Tspr4_3_V_1>>32'sd51)))) 
                  case (xpc10)
                      13'sd482/*482:xpc10*/:  xpc10 <= 13'sd483/*483:xpc10*/;

                      13'sd575/*575:xpc10*/:  xpc10 <= 13'sd576/*576:xpc10*/;

                      13'sd669/*669:xpc10*/:  xpc10 <= 13'sd670/*670:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd482/*482:xpc10*/:  xpc10 <= 13'sd4381/*4381:xpc10*/;

                      13'sd575/*575:xpc10*/:  xpc10 <= 13'sd3812/*3812:xpc10*/;

                      13'sd669/*669:xpc10*/:  xpc10 <= 13'sd3190/*3190:xpc10*/;
                  endcase
              if ((32'sd4094/*4094:USA10*/==(64'shfff&(Tspr4_3_V_0>>32'sd51)))) 
                  case (xpc10)
                      13'sd472/*472:xpc10*/:  xpc10 <= 13'sd473/*473:xpc10*/;

                      13'sd565/*565:xpc10*/:  xpc10 <= 13'sd566/*566:xpc10*/;

                      13'sd659/*659:xpc10*/:  xpc10 <= 13'sd660/*660:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd472/*472:xpc10*/:  xpc10 <= 13'sd4385/*4385:xpc10*/;

                      13'sd565/*565:xpc10*/:  xpc10 <= 13'sd3816/*3816:xpc10*/;

                      13'sd659/*659:xpc10*/:  xpc10 <= 13'sd3194/*3194:xpc10*/;
                  endcase
              if ((Tsfl0_9_V_6==32'sd0/*0:Tsfl0.9_V_6*/)) 
                  case (xpc10)
                      13'sd458/*458:xpc10*/:  xpc10 <= 13'sd459/*459:xpc10*/;

                      13'sd4503/*4503:xpc10*/:  xpc10 <= 13'sd4504/*4504:xpc10*/;

                      13'sd4532/*4532:xpc10*/:  xpc10 <= 13'sd4533/*4533:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd458/*458:xpc10*/:  xpc10 <= 13'sd468/*468:xpc10*/;

                      13'sd4503/*4503:xpc10*/:  xpc10 <= 13'sd4510/*4510:xpc10*/;

                      13'sd4532/*4532:xpc10*/:  xpc10 <= 13'sd4550/*4550:xpc10*/;
                  endcase
              if (!(!Tsfl0_9_V_3)) 
                  case (xpc10)
                      13'sd4499/*4499:xpc10*/:  xpc10 <= 13'sd4510/*4510:xpc10*/;

                      13'sd4528/*4528:xpc10*/:  xpc10 <= 13'sd4588/*4588:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd4499/*4499:xpc10*/:  xpc10 <= 13'sd4500/*4500:xpc10*/;

                      13'sd4528/*4528:xpc10*/:  xpc10 <= 13'sd4529/*4529:xpc10*/;
                  endcase
              if (!(!Tsfl0_9_V_4)) 
                  case (xpc10)
                      13'sd4391/*4391:xpc10*/:  xpc10 <= 13'sd4402/*4402:xpc10*/;

                      13'sd4590/*4590:xpc10*/:  xpc10 <= 13'sd4650/*4650:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd4391/*4391:xpc10*/:  xpc10 <= 13'sd4392/*4392:xpc10*/;

                      13'sd4590/*4590:xpc10*/:  xpc10 <= 13'sd4591/*4591:xpc10*/;
                  endcase
              if (!(!Tsfl1_8_V_3)) 
                  case (xpc10)
                      13'sd3930/*3930:xpc10*/:  xpc10 <= 13'sd3941/*3941:xpc10*/;

                      13'sd3959/*3959:xpc10*/:  xpc10 <= 13'sd4019/*4019:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd3930/*3930:xpc10*/:  xpc10 <= 13'sd3931/*3931:xpc10*/;

                      13'sd3959/*3959:xpc10*/:  xpc10 <= 13'sd3960/*3960:xpc10*/;
                  endcase
              if (!(!Tsfl1_8_V_4)) 
                  case (xpc10)
                      13'sd3822/*3822:xpc10*/:  xpc10 <= 13'sd3833/*3833:xpc10*/;

                      13'sd4021/*4021:xpc10*/:  xpc10 <= 13'sd4081/*4081:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd3822/*3822:xpc10*/:  xpc10 <= 13'sd3823/*3823:xpc10*/;

                      13'sd4021/*4021:xpc10*/:  xpc10 <= 13'sd4022/*4022:xpc10*/;
                  endcase
              if (Tsin1_19_V_0) 
                  case (xpc10)
                      13'sd3742/*3742:xpc10*/:  xpc10 <= 13'sd3743/*3743:xpc10*/;

                      13'sd3774/*3774:xpc10*/:  xpc10 <= 13'sd3775/*3775:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd3742/*3742:xpc10*/:  xpc10 <= 13'sd3788/*3788:xpc10*/;

                      13'sd3774/*3774:xpc10*/:  xpc10 <= 13'sd3784/*3784:xpc10*/;
                  endcase
              if (!(!Tsfl1_24_V_3)) 
                  case (xpc10)
                      13'sd3308/*3308:xpc10*/:  xpc10 <= 13'sd3319/*3319:xpc10*/;

                      13'sd3337/*3337:xpc10*/:  xpc10 <= 13'sd3397/*3397:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd3308/*3308:xpc10*/:  xpc10 <= 13'sd3309/*3309:xpc10*/;

                      13'sd3337/*3337:xpc10*/:  xpc10 <= 13'sd3338/*3338:xpc10*/;
                  endcase
              if (!(!Tsfl1_24_V_4)) 
                  case (xpc10)
                      13'sd3200/*3200:xpc10*/:  xpc10 <= 13'sd3211/*3211:xpc10*/;

                      13'sd3399/*3399:xpc10*/:  xpc10 <= 13'sd3459/*3459:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd3200/*3200:xpc10*/:  xpc10 <= 13'sd3201/*3201:xpc10*/;

                      13'sd3399/*3399:xpc10*/:  xpc10 <= 13'sd3400/*3400:xpc10*/;
                  endcase
              if ((Tsco5_4_V_0<32'sh100_0000)) 
                  case (xpc10)
                      13'sd3140/*3140:xpc10*/:  xpc10 <= 13'sd3141/*3141:xpc10*/;

                      13'sd3762/*3762:xpc10*/:  xpc10 <= 13'sd3763/*3763:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd3140/*3140:xpc10*/:  xpc10 <= 13'sd3147/*3147:xpc10*/;

                      13'sd3762/*3762:xpc10*/:  xpc10 <= 13'sd3769/*3769:xpc10*/;
                  endcase
              if ((Tsco5_4_V_0<32'sh1_0000)) 
                  case (xpc10)
                      13'sd3131/*3131:xpc10*/:  xpc10 <= 13'sd3132/*3132:xpc10*/;

                      13'sd3753/*3753:xpc10*/:  xpc10 <= 13'sd3754/*3754:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd3131/*3131:xpc10*/:  xpc10 <= 13'sd3138/*3138:xpc10*/;

                      13'sd3753/*3753:xpc10*/:  xpc10 <= 13'sd3760/*3760:xpc10*/;
                  endcase
              if (Tsin1_34_V_0) 
                  case (xpc10)
                      13'sd3120/*3120:xpc10*/:  xpc10 <= 13'sd3121/*3121:xpc10*/;

                      13'sd3152/*3152:xpc10*/:  xpc10 <= 13'sd3153/*3153:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd3120/*3120:xpc10*/:  xpc10 <= 13'sd3166/*3166:xpc10*/;

                      13'sd3152/*3152:xpc10*/:  xpc10 <= 13'sd3162/*3162:xpc10*/;
                  endcase
              if ((Tsmu5_7_V_5<Tsmu5_7_V_6)) 
                  case (xpc10)
                      13'sd2972/*2972:xpc10*/:  xpc10 <= 13'sd2973/*2973:xpc10*/;

                      13'sd2984/*2984:xpc10*/:  xpc10 <= 13'sd2985/*2985:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd2972/*2972:xpc10*/:  xpc10 <= 13'sd3093/*3093:xpc10*/;

                      13'sd2984/*2984:xpc10*/:  xpc10 <= 13'sd3088/*3088:xpc10*/;
                  endcase
              if ((Tsro33_4_V_1==32'sd0/*0:Tsro33.4_V_1*/)) 
                  case (xpc10)
                      13'sd2840/*2840:xpc10*/:  xpc10 <= 13'sd2841/*2841:xpc10*/;

                      13'sd2889/*2889:xpc10*/:  xpc10 <= 13'sd2899/*2899:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd2840/*2840:xpc10*/:  xpc10 <= 13'sd2846/*2846:xpc10*/;

                      13'sd2889/*2889:xpc10*/:  xpc10 <= 13'sd2890/*2890:xpc10*/;
                  endcase
              if (!(!Tsro33_4_V_6)) 
                  case (xpc10)
                      13'sd2815/*2815:xpc10*/:  xpc10 <= 13'sd2816/*2816:xpc10*/;

                      13'sd2823/*2823:xpc10*/:  xpc10 <= 13'sd2824/*2824:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd2815/*2815:xpc10*/:  xpc10 <= 13'sd2821/*2821:xpc10*/;

                      13'sd2823/*2823:xpc10*/:  xpc10 <= 13'sd2829/*2829:xpc10*/;
                  endcase
              if ((Tsmu26_4_V_5<Tsmu26_4_V_6)) 
                  case (xpc10)
                      13'sd2657/*2657:xpc10*/:  xpc10 <= 13'sd2658/*2658:xpc10*/;

                      13'sd2669/*2669:xpc10*/:  xpc10 <= 13'sd2670/*2670:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd2657/*2657:xpc10*/:  xpc10 <= 13'sd2947/*2947:xpc10*/;

                      13'sd2669/*2669:xpc10*/:  xpc10 <= 13'sd2942/*2942:xpc10*/;
                  endcase
              if (!(!Tsfl1_35_V_3)) 
                  case (xpc10)
                      13'sd2493/*2493:xpc10*/:  xpc10 <= 13'sd2504/*2504:xpc10*/;

                      13'sd2561/*2561:xpc10*/:  xpc10 <= 13'sd2621/*2621:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd2493/*2493:xpc10*/:  xpc10 <= 13'sd2494/*2494:xpc10*/;

                      13'sd2561/*2561:xpc10*/:  xpc10 <= 13'sd2562/*2562:xpc10*/;
                  endcase
              if ((Tsfl1_35_V_4==32'sd2047/*2047:Tsfl1.35_V_4*/)) 
                  case (xpc10)
                      13'sd2290/*2290:xpc10*/:  xpc10 <= 13'sd2291/*2291:xpc10*/;

                      13'sd2390/*2390:xpc10*/:  xpc10 <= 13'sd2391/*2391:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd2290/*2290:xpc10*/:  xpc10 <= 13'sd2372/*2372:xpc10*/;

                      13'sd2390/*2390:xpc10*/:  xpc10 <= 13'sd2483/*2483:xpc10*/;
                  endcase
              if (!(!Tssu2_4_V_1)) 
                  case (xpc10)
                      13'sd2062/*2062:xpc10*/:  xpc10 <= 13'sd2128/*2128:xpc10*/;

                      13'sd2222/*2222:xpc10*/:  xpc10 <= 13'sd2229/*2229:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd2062/*2062:xpc10*/:  xpc10 <= 13'sd2063/*2063:xpc10*/;

                      13'sd2222/*2222:xpc10*/:  xpc10 <= 13'sd2223/*2223:xpc10*/;
                  endcase
              if ((Tsro0_16_V_1==32'sd0/*0:Tsro0.16_V_1*/)) 
                  case (xpc10)
                      13'sd1846/*1846:xpc10*/:  xpc10 <= 13'sd1847/*1847:xpc10*/;

                      13'sd1895/*1895:xpc10*/:  xpc10 <= 13'sd1905/*1905:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd1846/*1846:xpc10*/:  xpc10 <= 13'sd1852/*1852:xpc10*/;

                      13'sd1895/*1895:xpc10*/:  xpc10 <= 13'sd1896/*1896:xpc10*/;
                  endcase
              if (!(!Tsro0_16_V_6)) 
                  case (xpc10)
                      13'sd1821/*1821:xpc10*/:  xpc10 <= 13'sd1822/*1822:xpc10*/;

                      13'sd1829/*1829:xpc10*/:  xpc10 <= 13'sd1830/*1830:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd1821/*1821:xpc10*/:  xpc10 <= 13'sd1827/*1827:xpc10*/;

                      13'sd1829/*1829:xpc10*/:  xpc10 <= 13'sd1835/*1835:xpc10*/;
                  endcase
              if (Tssu2_4_V_0) 
                  case (xpc10)
                      13'sd1765/*1765:xpc10*/:  xpc10 <= 13'sd1766/*1766:xpc10*/;

                      13'sd1854/*1854:xpc10*/:  xpc10 <= 13'sd1855/*1855:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd1765/*1765:xpc10*/:  xpc10 <= 13'sd1796/*1796:xpc10*/;

                      13'sd1854/*1854:xpc10*/:  xpc10 <= 13'sd1864/*1864:xpc10*/;
                  endcase
              if ((Tssu2_4_V_1==32'sd2047/*2047:Tssu2.4_V_1*/)) 
                  case (xpc10)
                      13'sd1592/*1592:xpc10*/:  xpc10 <= 13'sd1593/*1593:xpc10*/;

                      13'sd2134/*2134:xpc10*/:  xpc10 <= 13'sd2135/*2135:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd1592/*1592:xpc10*/:  xpc10 <= 13'sd1677/*1677:xpc10*/;

                      13'sd2134/*2134:xpc10*/:  xpc10 <= 13'sd2220/*2220:xpc10*/;
                  endcase
              if (!(!Tsad1_3_V_0)) 
                  case (xpc10)
                      13'sd1399/*1399:xpc10*/:  xpc10 <= 13'sd1459/*1459:xpc10*/;

                      13'sd1552/*1552:xpc10*/:  xpc10 <= 13'sd1570/*1570:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd1399/*1399:xpc10*/:  xpc10 <= 13'sd1400/*1400:xpc10*/;

                      13'sd1552/*1552:xpc10*/:  xpc10 <= 13'sd1553/*1553:xpc10*/;
                  endcase
              if ((Tsro28_4_V_1==32'sd0/*0:Tsro28.4_V_1*/)) 
                  case (xpc10)
                      13'sd1190/*1190:xpc10*/:  xpc10 <= 13'sd1191/*1191:xpc10*/;

                      13'sd1239/*1239:xpc10*/:  xpc10 <= 13'sd1249/*1249:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd1190/*1190:xpc10*/:  xpc10 <= 13'sd1196/*1196:xpc10*/;

                      13'sd1239/*1239:xpc10*/:  xpc10 <= 13'sd1240/*1240:xpc10*/;
                  endcase
              if (!(!Tsro28_4_V_6)) 
                  case (xpc10)
                      13'sd1165/*1165:xpc10*/:  xpc10 <= 13'sd1166/*1166:xpc10*/;

                      13'sd1173/*1173:xpc10*/:  xpc10 <= 13'sd1174/*1174:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd1165/*1165:xpc10*/:  xpc10 <= 13'sd1171/*1171:xpc10*/;

                      13'sd1173/*1173:xpc10*/:  xpc10 <= 13'sd1179/*1179:xpc10*/;
                  endcase
              if ((Tsad1_3_V_0==32'sd2047/*2047:Tsad1.3_V_0*/)) 
                  case (xpc10)
                      13'sd816/*816:xpc10*/:  xpc10 <= 13'sd817/*817:xpc10*/;

                      13'sd1465/*1465:xpc10*/:  xpc10 <= 13'sd1466/*1466:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd816/*816:xpc10*/:  xpc10 <= 13'sd1048/*1048:xpc10*/;

                      13'sd1465/*1465:xpc10*/:  xpc10 <= 13'sd1550/*1550:xpc10*/;
                  endcase
              if ((Tsfl1_24_V_4==32'sd2047/*2047:Tsfl1.24_V_4*/)) 
                  case (xpc10)
                      13'sd649/*649:xpc10*/:  xpc10 <= 13'sd650/*650:xpc10*/;

                      13'sd3229/*3229:xpc10*/:  xpc10 <= 13'sd3230/*3230:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd649/*649:xpc10*/:  xpc10 <= 13'sd3198/*3198:xpc10*/;

                      13'sd3229/*3229:xpc10*/:  xpc10 <= 13'sd3335/*3335:xpc10*/;
                  endcase
              if (!(!(32'sd2*Tdsi1_5_V_2*(32'sd1+32'sd2*Tdsi1_5_V_2)))) 
                  case (xpc10)
                      13'sd606/*606:xpc10*/:  xpc10 <= 13'sd3739/*3739:xpc10*/;

                      13'sd700/*700:xpc10*/:  xpc10 <= 13'sd3117/*3117:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd606/*606:xpc10*/:  xpc10 <= 13'sd607/*607:xpc10*/;

                      13'sd700/*700:xpc10*/:  xpc10 <= 13'sd701/*701:xpc10*/;
                  endcase
              if ((Tsfl1_8_V_4==32'sd2047/*2047:Tsfl1.8_V_4*/)) 
                  case (xpc10)
                      13'sd555/*555:xpc10*/:  xpc10 <= 13'sd556/*556:xpc10*/;

                      13'sd3851/*3851:xpc10*/:  xpc10 <= 13'sd3852/*3852:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd555/*555:xpc10*/:  xpc10 <= 13'sd3820/*3820:xpc10*/;

                      13'sd3851/*3851:xpc10*/:  xpc10 <= 13'sd3957/*3957:xpc10*/;
                  endcase
              if ((64'sh0<(Tdsi1_5_V_3>>32'sd63))) 
                  case (xpc10)
                      13'sd537/*537:xpc10*/:  xpc10 <= 13'sd538/*538:xpc10*/;

                      13'sd631/*631:xpc10*/:  xpc10 <= 13'sd632/*632:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd537/*537:xpc10*/:  xpc10 <= 13'sd4353/*4353:xpc10*/;

                      13'sd631/*631:xpc10*/:  xpc10 <= 13'sd3731/*3731:xpc10*/;
                  endcase
              if ((Tsfl0_9_V_4==32'sd2047/*2047:Tsfl0.9_V_4*/)) 
                  case (xpc10)
                      13'sd462/*462:xpc10*/:  xpc10 <= 13'sd463/*463:xpc10*/;

                      13'sd4420/*4420:xpc10*/:  xpc10 <= 13'sd4421/*4421:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd462/*462:xpc10*/:  xpc10 <= 13'sd4389/*4389:xpc10*/;

                      13'sd4420/*4420:xpc10*/:  xpc10 <= 13'sd4526/*4526:xpc10*/;
                  endcase
              if ((64'sh0<(A_64_US_CC_SCALbx12_ARB0[Tdbm0_3_V_1]>>32'sd63))) 
                  case (xpc10)
                      13'sd433/*433:xpc10*/:  xpc10 <= 13'sd434/*434:xpc10*/;

                      13'sd444/*444:xpc10*/:  xpc10 <= 13'sd445/*445:xpc10*/;
                  endcase
                   else 
                  case (xpc10)
                      13'sd433/*433:xpc10*/:  xpc10 <= 13'sd4926/*4926:xpc10*/;

                      13'sd444/*444:xpc10*/:  xpc10 <= 13'sd4922/*4922:xpc10*/;
                  endcase
              if (!Tspr11_2_V_2 && !Tspr11_2_V_4) 
                  case (xpc10)
                      13'sd3260/*3260:xpc10*/:  xpc10 <= 13'sd3266/*3266:xpc10*/;

                      13'sd3882/*3882:xpc10*/:  xpc10 <= 13'sd3888/*3888:xpc10*/;

                      13'sd4451/*4451:xpc10*/:  xpc10 <= 13'sd4457/*4457:xpc10*/;
                  endcase
                  if (Tspr11_2_V_2 || Tspr11_2_V_4) 
                  case (xpc10)
                      13'sd3260/*3260:xpc10*/:  xpc10 <= 13'sd3261/*3261:xpc10*/;

                      13'sd3882/*3882:xpc10*/:  xpc10 <= 13'sd3883/*3883:xpc10*/;

                      13'sd4451/*4451:xpc10*/:  xpc10 <= 13'sd4452/*4452:xpc10*/;
                  endcase
                  if (!Tspr4_3_V_2 && !Tspr4_3_V_4) 
                  case (xpc10)
                      13'sd493/*493:xpc10*/:  xpc10 <= 13'sd499/*499:xpc10*/;

                      13'sd586/*586:xpc10*/:  xpc10 <= 13'sd592/*592:xpc10*/;

                      13'sd680/*680:xpc10*/:  xpc10 <= 13'sd686/*686:xpc10*/;
                  endcase
                  if (Tspr4_3_V_2 || Tspr4_3_V_4) 
                  case (xpc10)
                      13'sd493/*493:xpc10*/:  xpc10 <= 13'sd494/*494:xpc10*/;

                      13'sd586/*586:xpc10*/:  xpc10 <= 13'sd587/*587:xpc10*/;

                      13'sd680/*680:xpc10*/:  xpc10 <= 13'sd681/*681:xpc10*/;
                  endcase
                  
              case (xpc10)
                  13'sd4710/*4710:xpc10*/:  begin 
                       xpc10 <= 13'sd4711/*4711:xpc10*/;
                       Tsf0_SPILL_259 <= 64'sh1;
                       end 
                      
                  13'sd4711/*4711:xpc10*/:  begin 
                       xpc10 <= 13'sd4712/*4712:xpc10*/;
                       Tsf0_SPILL_258 <= Tsf0_SPILL_257;
                       end 
                      
                  13'sd4715/*4715:xpc10*/:  begin 
                       xpc10 <= 13'sd4716/*4716:xpc10*/;
                       Tsfl0_9_V_8 <= Tsf0_SPILL_259|Tsf0_SPILL_258;
                       end 
                      
                  13'sd4716/*4716:xpc10*/: if (((Tsfl0_9_V_8<<32'sd1)<64'sh0))  xpc10 <= 13'sd4723/*4723:xpc10*/;
                       else  xpc10 <= 13'sd4717/*4717:xpc10*/;

                  13'sd4720/*4720:xpc10*/:  begin 
                       xpc10 <= 13'sd4721/*4721:xpc10*/;
                       Tsfl0_9_V_8 <= (Tsfl0_9_V_8<<32'sd1);
                       end 
                      
                  13'sd4721/*4721:xpc10*/:  begin 
                       xpc10 <= 13'sd4722/*4722:xpc10*/;
                       Tsfl0_9_V_5 <= rtl_signed_bitextract0(-16'sd1+Tsfl0_9_V_5);
                       end 
                      
                  13'sd4725/*4725:xpc10*/:  begin 
                       xpc10 <= 13'sd4726/*4726:xpc10*/;
                       Tsro29_4_V_0 <= rtl_signed_bitextract0(Tsfl0_9_V_5);
                       end 
                      
                  13'sd4726/*4726:xpc10*/:  begin 
                       xpc10 <= 13'sd4727/*4727:xpc10*/;
                       Tsro29_4_V_1 <= Tsfl0_9_V_8;
                       end 
                      
                  13'sd4729/*4729:xpc10*/:  begin 
                       xpc10 <= 13'sd4730/*4730:xpc10*/;
                       Tsro29_4_V_5 <= 16'sh200;
                       end 
                      
                  13'sd4733/*4733:xpc10*/:  begin 
                       xpc10 <= 13'sd4734/*4734:xpc10*/;
                       Tsro29_4_V_6 <= rtl_signed_bitextract2(64'sh3ff&Tsro29_4_V_1);
                       end 
                      
                  13'sd4755/*4755:xpc10*/:  begin 
                       xpc10 <= 13'sd4756/*4756:xpc10*/;
                       Tsp13_SPILL_256 <= 64'sh1;
                       end 
                      
                  13'sd4759/*4759:xpc10*/:  begin 
                       xpc10 <= 13'sd4760/*4760:xpc10*/;
                       fastspilldup24 <= $signed(64'sh_7ff0_0000_0000_0000+(Tsp13_SPILL_256<<32'sd63));
                       end 
                      
                  13'sd4760/*4760:xpc10*/:  begin 
                       xpc10 <= 13'sd4761/*4761:xpc10*/;
                       Tsr29_SPILL_260 <= fastspilldup24;
                       end 
                      
                  13'sd4761/*4761:xpc10*/:  begin 
                       xpc10 <= 13'sd4762/*4762:xpc10*/;
                       Tsr29_SPILL_256 <= fastspilldup24;
                       end 
                      
                  13'sd4766/*4766:xpc10*/:  begin 
                       xpc10 <= 13'sd4767/*4767:xpc10*/;
                       Tsr29_SPILL_258 <= 64'sh1;
                       end 
                      
                  13'sd4767/*4767:xpc10*/:  begin 
                       xpc10 <= 13'sd4768/*4768:xpc10*/;
                       Tsr29_SPILL_257 <= Tsr29_SPILL_256;
                       end 
                      
                  13'sd4771/*4771:xpc10*/:  begin 
                       xpc10 <= 13'sd4772/*4772:xpc10*/;
                       Tsr29_SPILL_259 <= Tsr29_SPILL_257+(0-Tsr29_SPILL_258);
                       end 
                      
                  13'sd4775/*4775:xpc10*/:  begin 
                       xpc10 <= 13'sd4776/*4776:xpc10*/;
                       Tsf0_SPILL_256 <= Tsr29_SPILL_259;
                       end 
                      
                  13'sd4779/*4779:xpc10*/:  begin 
                       xpc10 <= 13'sd4780/*4780:xpc10*/;
                       Tsr29_SPILL_258 <= 64'sh0;
                       end 
                      
                  13'sd4780/*4780:xpc10*/:  begin 
                       xpc10 <= 13'sd4781/*4781:xpc10*/;
                       Tsr29_SPILL_257 <= Tsr29_SPILL_260;
                       end 
                      
                  13'sd4784/*4784:xpc10*/:  begin 
                       xpc10 <= 13'sd4785/*4785:xpc10*/;
                       Tsp13_SPILL_256 <= 64'sh0;
                       end 
                      
                  13'sd4797/*4797:xpc10*/:  begin 
                       xpc10 <= 13'sd4798/*4798:xpc10*/;
                       Tssh18_7_V_0 <= Tsro29_4_V_1;
                       end 
                      
                  13'sd4801/*4801:xpc10*/:  begin 
                       xpc10 <= 13'sd4802/*4802:xpc10*/;
                       Tsro29_4_V_1 <= Tssh18_7_V_0;
                       end 
                      
                  13'sd4802/*4802:xpc10*/:  begin 
                       xpc10 <= 13'sd4803/*4803:xpc10*/;
                       Tsro29_4_V_0 <= 16'sh0;
                       end 
                      
                  13'sd4803/*4803:xpc10*/:  begin 
                       xpc10 <= 13'sd4804/*4804:xpc10*/;
                       Tsro29_4_V_6 <= rtl_signed_bitextract2(64'sh3ff&Tsro29_4_V_1);
                       end 
                      
                  13'sd4823/*4823:xpc10*/:  begin 
                       xpc10 <= 13'sd4824/*4824:xpc10*/;
                       Tsro29_4_V_1 <= (Tsro29_4_V_1+rtl_sign_extend1(Tsro29_4_V_5)>>32'sd10);
                       end 
                      
                  13'sd4828/*4828:xpc10*/:  begin 
                       xpc10 <= 13'sd4829/*4829:xpc10*/;
                       Tsro29_4_V_1 <= -64'sh2&Tsro29_4_V_1;
                       end 
                      
                  13'sd4836/*4836:xpc10*/:  begin 
                       xpc10 <= 13'sd4837/*4837:xpc10*/;
                       Tsro29_4_V_0 <= 16'sh0;
                       end 
                      
                  13'sd4844/*4844:xpc10*/:  begin 
                       xpc10 <= 13'sd4845/*4845:xpc10*/;
                       Tsp27_SPILL_256 <= 64'sh1;
                       end 
                      
                  13'sd4848/*4848:xpc10*/:  begin 
                       xpc10 <= 13'sd4849/*4849:xpc10*/;
                       Tsr29_SPILL_259 <= Tsro29_4_V_1+(Tsp27_SPILL_256<<32'sd63)+(rtl_sign_extend1(Tsro29_4_V_0)<<32'sd52);
                       end 
                      
                  13'sd4852/*4852:xpc10*/:  begin 
                       xpc10 <= 13'sd4853/*4853:xpc10*/;
                       Tsp27_SPILL_256 <= 64'sh0;
                       end 
                      
                  13'sd4860/*4860:xpc10*/:  begin 
                       xpc10 <= 13'sd4861/*4861:xpc10*/;
                       fastspilldup26 <= (Tsro29_4_V_1>>(32'sd63&rtl_signed_bitextract0((0-Tsro29_4_V_0))));
                       end 
                      
                  13'sd4861/*4861:xpc10*/:  begin 
                       xpc10 <= 13'sd4862/*4862:xpc10*/;
                       Tss18_SPILL_259 <= fastspilldup26;
                       end 
                      
                  13'sd4862/*4862:xpc10*/:  begin 
                       xpc10 <= 13'sd4863/*4863:xpc10*/;
                       Tss18_SPILL_256 <= fastspilldup26;
                       end 
                      
                  13'sd4867/*4867:xpc10*/:  begin 
                       xpc10 <= 13'sd4868/*4868:xpc10*/;
                       Tss18_SPILL_258 <= 64'sh1;
                       end 
                      
                  13'sd4868/*4868:xpc10*/:  begin 
                       xpc10 <= 13'sd4869/*4869:xpc10*/;
                       Tss18_SPILL_257 <= Tss18_SPILL_256;
                       end 
                      
                  13'sd4872/*4872:xpc10*/:  begin 
                       xpc10 <= 13'sd4873/*4873:xpc10*/;
                       Tssh18_7_V_0 <= Tss18_SPILL_258|Tss18_SPILL_257;
                       end 
                      
                  13'sd4876/*4876:xpc10*/:  begin 
                       xpc10 <= 13'sd4877/*4877:xpc10*/;
                       Tss18_SPILL_258 <= 64'sh0;
                       end 
                      
                  13'sd4877/*4877:xpc10*/:  begin 
                       xpc10 <= 13'sd4878/*4878:xpc10*/;
                       Tss18_SPILL_257 <= Tss18_SPILL_259;
                       end 
                      
                  13'sd4885/*4885:xpc10*/:  begin 
                       xpc10 <= 13'sd4886/*4886:xpc10*/;
                       Tss18_SPILL_260 <= 64'sh1;
                       end 
                      
                  13'sd4889/*4889:xpc10*/:  begin 
                       xpc10 <= 13'sd4890/*4890:xpc10*/;
                       Tssh18_7_V_0 <= Tss18_SPILL_260;
                       end 
                      
                  13'sd4893/*4893:xpc10*/:  begin 
                       xpc10 <= 13'sd4894/*4894:xpc10*/;
                       Tss18_SPILL_260 <= 64'sh0;
                       end 
                      
                  13'sd4897/*4897:xpc10*/:  begin 
                       xpc10 <= 13'sd4898/*4898:xpc10*/;
                       Tsf0_SPILL_259 <= 64'sh0;
                       end 
                      
                  13'sd4898/*4898:xpc10*/:  begin 
                       xpc10 <= 13'sd4899/*4899:xpc10*/;
                       Tsf0_SPILL_258 <= Tsf0_SPILL_260;
                       end 
                      
                  13'sd4902/*4902:xpc10*/:  begin 
                       xpc10 <= 13'sd4903/*4903:xpc10*/;
                       Tsm24_SPILL_262 <= 64'sh0;
                       end 
                      
                  13'sd4903/*4903:xpc10*/:  begin 
                       xpc10 <= 13'sd4904/*4904:xpc10*/;
                       Tsm24_SPILL_261 <= Tsm24_SPILL_263;
                       end 
                      
                  13'sd4907/*4907:xpc10*/:  begin 
                       xpc10 <= 13'sd4908/*4908:xpc10*/;
                       Tsm24_SPILL_259 <= 64'sh0;
                       end 
                      
                  13'sd4908/*4908:xpc10*/:  begin 
                       xpc10 <= 13'sd4909/*4909:xpc10*/;
                       Tsm24_SPILL_258 <= Tsm24_SPILL_264;
                       end 
                      
                  13'sd4916/*4916:xpc10*/:  begin 
                       xpc10 <= 13'sd4917/*4917:xpc10*/;
                       Tsco0_2_V_0 <= (Tsco0_2_V_0>>32'sd32);
                       end 
                      
                  13'sd4920/*4920:xpc10*/:  begin 
                       xpc10 <= 13'sd4921/*4921:xpc10*/;
                       Tsco0_2_V_0 <= (Tsco0_2_V_0>>32'sd32);
                       end 
                      
                  13'sd4924/*4924:xpc10*/:  begin 
                       xpc10 <= 13'sd4925/*4925:xpc10*/;
                       Tse0SPILL10_256 <= 32'sd0;
                       end 
                      
                  13'sd4928/*4928:xpc10*/:  begin 
                       xpc10 <= 13'sd4929/*4929:xpc10*/;
                       Tse0_SPILL_256 <= 32'sd0;
                       end 
                      endcase
              if ((Tsfl0_9_V_9==32'sd0/*0:Tsfl0.9_V_9*/))  begin if ((13'sd4706/*4706:xpc10*/==xpc10))  xpc10 <= 13'sd4895/*4895:xpc10*/;
                       end 
                   else if ((13'sd4706/*4706:xpc10*/==xpc10))  xpc10 <= 13'sd4707/*4707:xpc10*/;
                      
              case (xpc10)
                  13'sd4141/*4141:xpc10*/:  begin 
                       xpc10 <= 13'sd4142/*4142:xpc10*/;
                       Tsf1_SPILL_259 <= 64'sh1;
                       end 
                      
                  13'sd4142/*4142:xpc10*/:  begin 
                       xpc10 <= 13'sd4143/*4143:xpc10*/;
                       Tsf1_SPILL_258 <= Tsf1_SPILL_257;
                       end 
                      
                  13'sd4146/*4146:xpc10*/:  begin 
                       xpc10 <= 13'sd4147/*4147:xpc10*/;
                       Tsfl1_8_V_8 <= Tsf1_SPILL_259|Tsf1_SPILL_258;
                       end 
                      
                  13'sd4147/*4147:xpc10*/: if (((Tsfl1_8_V_8<<32'sd1)<64'sh0))  xpc10 <= 13'sd4154/*4154:xpc10*/;
                       else  xpc10 <= 13'sd4148/*4148:xpc10*/;

                  13'sd4151/*4151:xpc10*/:  begin 
                       xpc10 <= 13'sd4152/*4152:xpc10*/;
                       Tsfl1_8_V_8 <= (Tsfl1_8_V_8<<32'sd1);
                       end 
                      
                  13'sd4152/*4152:xpc10*/:  begin 
                       xpc10 <= 13'sd4153/*4153:xpc10*/;
                       Tsfl1_8_V_5 <= rtl_signed_bitextract0(-16'sd1+Tsfl1_8_V_5);
                       end 
                      
                  13'sd4156/*4156:xpc10*/:  begin 
                       xpc10 <= 13'sd4157/*4157:xpc10*/;
                       Tsro29_4_V_0 <= rtl_signed_bitextract0(Tsfl1_8_V_5);
                       end 
                      
                  13'sd4157/*4157:xpc10*/:  begin 
                       xpc10 <= 13'sd4158/*4158:xpc10*/;
                       Tsro29_4_V_1 <= Tsfl1_8_V_8;
                       end 
                      
                  13'sd4160/*4160:xpc10*/:  begin 
                       xpc10 <= 13'sd4161/*4161:xpc10*/;
                       Tsro29_4_V_5 <= 16'sh200;
                       end 
                      
                  13'sd4164/*4164:xpc10*/:  begin 
                       xpc10 <= 13'sd4165/*4165:xpc10*/;
                       Tsro29_4_V_6 <= rtl_signed_bitextract2(64'sh3ff&Tsro29_4_V_1);
                       end 
                      
                  13'sd4186/*4186:xpc10*/:  begin 
                       xpc10 <= 13'sd4187/*4187:xpc10*/;
                       Tsp13_SPILL_256 <= 64'sh1;
                       end 
                      
                  13'sd4190/*4190:xpc10*/:  begin 
                       xpc10 <= 13'sd4191/*4191:xpc10*/;
                       fastspilldup34 <= $signed(64'sh_7ff0_0000_0000_0000+(Tsp13_SPILL_256<<32'sd63));
                       end 
                      
                  13'sd4191/*4191:xpc10*/:  begin 
                       xpc10 <= 13'sd4192/*4192:xpc10*/;
                       Tsr29_SPILL_260 <= fastspilldup34;
                       end 
                      
                  13'sd4192/*4192:xpc10*/:  begin 
                       xpc10 <= 13'sd4193/*4193:xpc10*/;
                       Tsr29_SPILL_256 <= fastspilldup34;
                       end 
                      
                  13'sd4197/*4197:xpc10*/:  begin 
                       xpc10 <= 13'sd4198/*4198:xpc10*/;
                       Tsr29_SPILL_258 <= 64'sh1;
                       end 
                      
                  13'sd4198/*4198:xpc10*/:  begin 
                       xpc10 <= 13'sd4199/*4199:xpc10*/;
                       Tsr29_SPILL_257 <= Tsr29_SPILL_256;
                       end 
                      
                  13'sd4202/*4202:xpc10*/:  begin 
                       xpc10 <= 13'sd4203/*4203:xpc10*/;
                       Tsr29_SPILL_259 <= Tsr29_SPILL_257+(0-Tsr29_SPILL_258);
                       end 
                      
                  13'sd4206/*4206:xpc10*/:  begin 
                       xpc10 <= 13'sd4207/*4207:xpc10*/;
                       Tsf1_SPILL_256 <= Tsr29_SPILL_259;
                       end 
                      
                  13'sd4210/*4210:xpc10*/:  begin 
                       xpc10 <= 13'sd4211/*4211:xpc10*/;
                       Tsr29_SPILL_258 <= 64'sh0;
                       end 
                      
                  13'sd4211/*4211:xpc10*/:  begin 
                       xpc10 <= 13'sd4212/*4212:xpc10*/;
                       Tsr29_SPILL_257 <= Tsr29_SPILL_260;
                       end 
                      
                  13'sd4215/*4215:xpc10*/:  begin 
                       xpc10 <= 13'sd4216/*4216:xpc10*/;
                       Tsp13_SPILL_256 <= 64'sh0;
                       end 
                      
                  13'sd4228/*4228:xpc10*/:  begin 
                       xpc10 <= 13'sd4229/*4229:xpc10*/;
                       Tssh18_7_V_0 <= Tsro29_4_V_1;
                       end 
                      
                  13'sd4232/*4232:xpc10*/:  begin 
                       xpc10 <= 13'sd4233/*4233:xpc10*/;
                       Tsro29_4_V_1 <= Tssh18_7_V_0;
                       end 
                      
                  13'sd4233/*4233:xpc10*/:  begin 
                       xpc10 <= 13'sd4234/*4234:xpc10*/;
                       Tsro29_4_V_0 <= 16'sh0;
                       end 
                      
                  13'sd4234/*4234:xpc10*/:  begin 
                       xpc10 <= 13'sd4235/*4235:xpc10*/;
                       Tsro29_4_V_6 <= rtl_signed_bitextract2(64'sh3ff&Tsro29_4_V_1);
                       end 
                      
                  13'sd4254/*4254:xpc10*/:  begin 
                       xpc10 <= 13'sd4255/*4255:xpc10*/;
                       Tsro29_4_V_1 <= (Tsro29_4_V_1+rtl_sign_extend1(Tsro29_4_V_5)>>32'sd10);
                       end 
                      
                  13'sd4259/*4259:xpc10*/:  begin 
                       xpc10 <= 13'sd4260/*4260:xpc10*/;
                       Tsro29_4_V_1 <= -64'sh2&Tsro29_4_V_1;
                       end 
                      
                  13'sd4267/*4267:xpc10*/:  begin 
                       xpc10 <= 13'sd4268/*4268:xpc10*/;
                       Tsro29_4_V_0 <= 16'sh0;
                       end 
                      
                  13'sd4275/*4275:xpc10*/:  begin 
                       xpc10 <= 13'sd4276/*4276:xpc10*/;
                       Tsp27_SPILL_256 <= 64'sh1;
                       end 
                      
                  13'sd4279/*4279:xpc10*/:  begin 
                       xpc10 <= 13'sd4280/*4280:xpc10*/;
                       Tsr29_SPILL_259 <= Tsro29_4_V_1+(Tsp27_SPILL_256<<32'sd63)+(rtl_sign_extend1(Tsro29_4_V_0)<<32'sd52);
                       end 
                      
                  13'sd4283/*4283:xpc10*/:  begin 
                       xpc10 <= 13'sd4284/*4284:xpc10*/;
                       Tsp27_SPILL_256 <= 64'sh0;
                       end 
                      
                  13'sd4291/*4291:xpc10*/:  begin 
                       xpc10 <= 13'sd4292/*4292:xpc10*/;
                       fastspilldup36 <= (Tsro29_4_V_1>>(32'sd63&rtl_signed_bitextract0((0-Tsro29_4_V_0))));
                       end 
                      
                  13'sd4292/*4292:xpc10*/:  begin 
                       xpc10 <= 13'sd4293/*4293:xpc10*/;
                       Tss18_SPILL_259 <= fastspilldup36;
                       end 
                      
                  13'sd4293/*4293:xpc10*/:  begin 
                       xpc10 <= 13'sd4294/*4294:xpc10*/;
                       Tss18_SPILL_256 <= fastspilldup36;
                       end 
                      
                  13'sd4298/*4298:xpc10*/:  begin 
                       xpc10 <= 13'sd4299/*4299:xpc10*/;
                       Tss18_SPILL_258 <= 64'sh1;
                       end 
                      
                  13'sd4299/*4299:xpc10*/:  begin 
                       xpc10 <= 13'sd4300/*4300:xpc10*/;
                       Tss18_SPILL_257 <= Tss18_SPILL_256;
                       end 
                      
                  13'sd4303/*4303:xpc10*/:  begin 
                       xpc10 <= 13'sd4304/*4304:xpc10*/;
                       Tssh18_7_V_0 <= Tss18_SPILL_258|Tss18_SPILL_257;
                       end 
                      
                  13'sd4307/*4307:xpc10*/:  begin 
                       xpc10 <= 13'sd4308/*4308:xpc10*/;
                       Tss18_SPILL_258 <= 64'sh0;
                       end 
                      
                  13'sd4308/*4308:xpc10*/:  begin 
                       xpc10 <= 13'sd4309/*4309:xpc10*/;
                       Tss18_SPILL_257 <= Tss18_SPILL_259;
                       end 
                      
                  13'sd4316/*4316:xpc10*/:  begin 
                       xpc10 <= 13'sd4317/*4317:xpc10*/;
                       Tss18_SPILL_260 <= 64'sh1;
                       end 
                      
                  13'sd4320/*4320:xpc10*/:  begin 
                       xpc10 <= 13'sd4321/*4321:xpc10*/;
                       Tssh18_7_V_0 <= Tss18_SPILL_260;
                       end 
                      
                  13'sd4324/*4324:xpc10*/:  begin 
                       xpc10 <= 13'sd4325/*4325:xpc10*/;
                       Tss18_SPILL_260 <= 64'sh0;
                       end 
                      
                  13'sd4328/*4328:xpc10*/:  begin 
                       xpc10 <= 13'sd4329/*4329:xpc10*/;
                       Tsf1_SPILL_259 <= 64'sh0;
                       end 
                      
                  13'sd4329/*4329:xpc10*/:  begin 
                       xpc10 <= 13'sd4330/*4330:xpc10*/;
                       Tsf1_SPILL_258 <= Tsf1_SPILL_260;
                       end 
                      
                  13'sd4333/*4333:xpc10*/:  begin 
                       xpc10 <= 13'sd4334/*4334:xpc10*/;
                       Tsm24_SPILL_262 <= 64'sh0;
                       end 
                      
                  13'sd4334/*4334:xpc10*/:  begin 
                       xpc10 <= 13'sd4335/*4335:xpc10*/;
                       Tsm24_SPILL_261 <= Tsm24_SPILL_263;
                       end 
                      
                  13'sd4338/*4338:xpc10*/:  begin 
                       xpc10 <= 13'sd4339/*4339:xpc10*/;
                       Tsm24_SPILL_259 <= 64'sh0;
                       end 
                      
                  13'sd4339/*4339:xpc10*/:  begin 
                       xpc10 <= 13'sd4340/*4340:xpc10*/;
                       Tsm24_SPILL_258 <= Tsm24_SPILL_264;
                       end 
                      
                  13'sd4347/*4347:xpc10*/:  begin 
                       xpc10 <= 13'sd4348/*4348:xpc10*/;
                       Tsco0_2_V_0 <= (Tsco0_2_V_0>>32'sd32);
                       end 
                      
                  13'sd4351/*4351:xpc10*/:  begin 
                       xpc10 <= 13'sd4352/*4352:xpc10*/;
                       Tsco0_2_V_0 <= (Tsco0_2_V_0>>32'sd32);
                       end 
                      
                  13'sd4355/*4355:xpc10*/:  begin 
                       xpc10 <= 13'sd4356/*4356:xpc10*/;
                       Tse0SPILL10_256 <= 32'sd0;
                       end 
                      
                  13'sd4359/*4359:xpc10*/:  begin 
                       xpc10 <= 13'sd4360/*4360:xpc10*/;
                       Tse0_SPILL_256 <= 32'sd0;
                       end 
                      
                  13'sd4367/*4367:xpc10*/:  begin 
                       xpc10 <= 13'sd4368/*4368:xpc10*/;
                       Tsp4_SPILL_256 <= Tspr4_3_V_0;
                       end 
                      
                  13'sd4375/*4375:xpc10*/:  begin 
                       xpc10 <= 13'sd4376/*4376:xpc10*/;
                       Tsp4_SPILL_256 <= Tspr4_3_V_1;
                       end 
                      
                  13'sd4379/*4379:xpc10*/:  begin 
                       xpc10 <= 13'sd4380/*4380:xpc10*/;
                       Tsp4_SPILL_256 <= Tspr4_3_V_0;
                       end 
                      
                  13'sd4383/*4383:xpc10*/:  begin 
                       xpc10 <= 13'sd4384/*4384:xpc10*/;
                       Tsf0SPILL12_256 <= 32'sd0;
                       end 
                      
                  13'sd4387/*4387:xpc10*/:  begin 
                       xpc10 <= 13'sd4388/*4388:xpc10*/;
                       Tsf0SPILL10_256 <= 32'sd0;
                       end 
                      
                  13'sd4400/*4400:xpc10*/:  begin 
                       xpc10 <= 13'sd4401/*4401:xpc10*/;
                       Tsf0_SPILL_256 <= 64'h_7fff_ffff_ffff_ffff;
                       end 
                      
                  13'sd4408/*4408:xpc10*/:  begin 
                       xpc10 <= 13'sd4409/*4409:xpc10*/;
                       Tsp8_SPILL_256 <= 64'sh1;
                       end 
                      
                  13'sd4412/*4412:xpc10*/:  begin 
                       xpc10 <= 13'sd4413/*4413:xpc10*/;
                       Tsf0_SPILL_256 <= $signed(64'sh_7ff0_0000_0000_0000+(Tsp8_SPILL_256<<32'sd63));
                       end 
                      
                  13'sd4416/*4416:xpc10*/:  begin 
                       xpc10 <= 13'sd4417/*4417:xpc10*/;
                       Tsp8_SPILL_256 <= 64'sh0;
                       end 
                      
                  13'sd4428/*4428:xpc10*/:  begin 
                       xpc10 <= 13'sd4429/*4429:xpc10*/;
                       Tspr11_2_V_0 <= $unsigned(A_64_US_CC_SCALbx12_ARB0[Tdbm0_3_V_1]);
                       end 
                      
                  13'sd4429/*4429:xpc10*/:  begin 
                       xpc10 <= 13'sd4430/*4430:xpc10*/;
                       Tspr11_2_V_1 <= $unsigned(A_64_US_CC_SCALbx12_ARB0[Tdbm0_3_V_1]);
                       end 
                      
                  13'sd4434/*4434:xpc10*/:  begin 
                       xpc10 <= 13'sd4435/*4435:xpc10*/;
                       Tsf0SPILL10_256 <= rtl_sign_extend3((32'sd0/*0:USA26*/==(32'sd0/*0:USA24*/==(64'sh7_ffff_ffff_ffff&Tspr11_2_V_0
                      ))));

                       end 
                      
                  13'sd4438/*4438:xpc10*/:  begin 
                       xpc10 <= 13'sd4439/*4439:xpc10*/;
                       Tspr11_2_V_2 <= rtl_unsigned_bitextract4(Tsf0SPILL10_256);
                       end 
                      
                  13'sd4439/*4439:xpc10*/:  begin 
                       xpc10 <= 13'sd4440/*4440:xpc10*/;
                       Tspr11_2_V_3 <= (32'sd0<rtl_sign_extend5(54'sd9007199254740992)+(Tspr11_2_V_1<<32'sd1));
                       end 
                      
                  13'sd4444/*4444:xpc10*/:  begin 
                       xpc10 <= 13'sd4445/*4445:xpc10*/;
                       Tsf0SPILL12_256 <= rtl_sign_extend3((32'sd0/*0:USA32*/==(32'sd0/*0:USA30*/==(64'sh7_ffff_ffff_ffff&Tspr11_2_V_1
                      ))));

                       end 
                      
                  13'sd4448/*4448:xpc10*/:  begin 
                       xpc10 <= 13'sd4449/*4449:xpc10*/;
                       Tspr11_2_V_4 <= rtl_unsigned_bitextract4(Tsf0SPILL12_256);
                       end 
                      
                  13'sd4449/*4449:xpc10*/:  begin 
                       xpc10 <= 13'sd4450/*4450:xpc10*/;
                       Tspr11_2_V_0 <= 64'sh8_0000_0000_0000|Tspr11_2_V_0;
                       end 
                      
                  13'sd4450/*4450:xpc10*/:  begin 
                       xpc10 <= 13'sd4451/*4451:xpc10*/;
                       Tspr11_2_V_1 <= 64'sh8_0000_0000_0000|Tspr11_2_V_1;
                       end 
                      
                  13'sd4463/*4463:xpc10*/:  begin 
                       xpc10 <= 13'sd4464/*4464:xpc10*/;
                       Tsp11_SPILL_256 <= Tspr11_2_V_1;
                       end 
                      
                  13'sd4467/*4467:xpc10*/:  begin 
                       xpc10 <= 13'sd4468/*4468:xpc10*/;
                       Tsf0_SPILL_256 <= Tsp11_SPILL_256;
                       end 
                      
                  13'sd4475/*4475:xpc10*/:  begin 
                       xpc10 <= 13'sd4476/*4476:xpc10*/;
                       Tsp11_SPILL_256 <= Tspr11_2_V_0;
                       end 
                      
                  13'sd4483/*4483:xpc10*/:  begin 
                       xpc10 <= 13'sd4484/*4484:xpc10*/;
                       Tsp11_SPILL_256 <= Tspr11_2_V_1;
                       end 
                      
                  13'sd4487/*4487:xpc10*/:  begin 
                       xpc10 <= 13'sd4488/*4488:xpc10*/;
                       Tsp11_SPILL_256 <= Tspr11_2_V_0;
                       end 
                      
                  13'sd4491/*4491:xpc10*/:  begin 
                       xpc10 <= 13'sd4492/*4492:xpc10*/;
                       Tsf0SPILL12_256 <= 32'sd0;
                       end 
                      
                  13'sd4495/*4495:xpc10*/:  begin 
                       xpc10 <= 13'sd4496/*4496:xpc10*/;
                       Tsf0SPILL10_256 <= 32'sd0;
                       end 
                      
                  13'sd4508/*4508:xpc10*/:  begin 
                       xpc10 <= 13'sd4509/*4509:xpc10*/;
                       Tsf0_SPILL_256 <= 64'h_7fff_ffff_ffff_ffff;
                       end 
                      
                  13'sd4516/*4516:xpc10*/:  begin 
                       xpc10 <= 13'sd4517/*4517:xpc10*/;
                       Tsp15_SPILL_256 <= 64'sh1;
                       end 
                      
                  13'sd4520/*4520:xpc10*/:  begin 
                       xpc10 <= 13'sd4521/*4521:xpc10*/;
                       Tsf0_SPILL_256 <= $signed(64'sh_7ff0_0000_0000_0000+(Tsp15_SPILL_256<<32'sd63));
                       end 
                      
                  13'sd4524/*4524:xpc10*/:  begin 
                       xpc10 <= 13'sd4525/*4525:xpc10*/;
                       Tsp15_SPILL_256 <= 64'sh0;
                       end 
                      
                  13'sd4540/*4540:xpc10*/:  begin 
                       xpc10 <= 13'sd4541/*4541:xpc10*/;
                       Tsp18_SPILL_256 <= 64'sh1;
                       end 
                      
                  13'sd4544/*4544:xpc10*/:  begin 
                       xpc10 <= 13'sd4545/*4545:xpc10*/;
                       Tsf0_SPILL_256 <= $signed(64'sh0+(Tsp18_SPILL_256<<32'sd63));
                       end 
                      
                  13'sd4548/*4548:xpc10*/:  begin 
                       xpc10 <= 13'sd4549/*4549:xpc10*/;
                       Tsp18_SPILL_256 <= 64'sh0;
                       end 
                      
                  13'sd4552/*4552:xpc10*/:  begin 
                       xpc10 <= 13'sd4553/*4553:xpc10*/;
                       Tsco0_2_V_0 <= Tsfl0_9_V_6;
                       end 
                      
                  13'sd4553/*4553:xpc10*/:  begin 
                       xpc10 <= 13'sd4554/*4554:xpc10*/;
                       Tsco0_2_V_1 <= 8'h0;
                       end 
                      
                  13'sd4558/*4558:xpc10*/:  begin 
                       xpc10 <= 13'sd4559/*4559:xpc10*/;
                       Tsco0_2_V_1 <= 8'h20;
                       end 
                      
                  13'sd4562/*4562:xpc10*/:  begin 
                       xpc10 <= 13'sd4563/*4563:xpc10*/;
                       Tsco3_7_V_0 <= rtl_unsigned_bitextract6(64'h_ffff_ffff&Tsco0_2_V_0);
                       end 
                      
                  13'sd4563/*4563:xpc10*/:  begin 
                       xpc10 <= 13'sd4564/*4564:xpc10*/;
                       Tsco3_7_V_1 <= 8'h0;
                       end 
                      
                  13'sd4568/*4568:xpc10*/:  begin 
                       xpc10 <= 13'sd4569/*4569:xpc10*/;
                       Tsco3_7_V_1 <= 8'h10;
                       end 
                      
                  13'sd4569/*4569:xpc10*/:  begin 
                       xpc10 <= 13'sd4570/*4570:xpc10*/;
                       Tsco3_7_V_0 <= (Tsco3_7_V_0<<32'sd16);
                       end 
                      
                  13'sd4577/*4577:xpc10*/:  begin 
                       xpc10 <= 13'sd4578/*4578:xpc10*/;
                       Tsco3_7_V_1 <= rtl_unsigned_bitextract7(8'd8+Tsco3_7_V_1);
                       end 
                      
                  13'sd4578/*4578:xpc10*/:  begin 
                       xpc10 <= 13'sd4579/*4579:xpc10*/;
                       Tsco3_7_V_0 <= (Tsco3_7_V_0<<32'sd8);
                       end 
                      
                  13'sd4582/*4582:xpc10*/:  begin 
                       xpc10 <= 13'sd4583/*4583:xpc10*/;
                       Tsco3_7_V_1 <= rtl_unsigned_bitextract7(Tsco3_7_V_1+A_8_US_CC_SCALbx16_ARA0[$unsigned((Tsco3_7_V_0>>32'sd24))]
                      );

                       end 
                      
                  13'sd4583/*4583:xpc10*/:  begin 
                       xpc10 <= 13'sd4584/*4584:xpc10*/;
                       Tsco0_2_V_1 <= rtl_unsigned_bitextract7(Tsco0_2_V_1+Tsco3_7_V_1);
                       end 
                      
                  13'sd4584/*4584:xpc10*/:  begin 
                       xpc10 <= 13'sd4585/*4585:xpc10*/;
                       Tsno19_4_V_0 <= $unsigned(-32'sd11+rtl_sign_extend8(Tsco0_2_V_1));
                       end 
                      
                  13'sd4585/*4585:xpc10*/:  begin 
                       xpc10 <= 13'sd4586/*4586:xpc10*/;
                       Tsfl0_9_V_6 <= (Tsfl0_9_V_6<<(32'sd63&Tsno19_4_V_0));
                       end 
                      
                  13'sd4586/*4586:xpc10*/:  begin 
                       xpc10 <= 13'sd4587/*4587:xpc10*/;
                       Tsfl0_9_V_3 <= rtl_signed_bitextract0(rtl_sign_extend9(16'sd1)+(0-Tsno19_4_V_0));
                       end 
                      
                  13'sd4602/*4602:xpc10*/:  begin 
                       xpc10 <= 13'sd4603/*4603:xpc10*/;
                       Tsp22_SPILL_256 <= 64'sh1;
                       end 
                      
                  13'sd4606/*4606:xpc10*/:  begin 
                       xpc10 <= 13'sd4607/*4607:xpc10*/;
                       Tsf0_SPILL_256 <= $signed(64'sh0+(Tsp22_SPILL_256<<32'sd63));
                       end 
                      
                  13'sd4610/*4610:xpc10*/:  begin 
                       xpc10 <= 13'sd4611/*4611:xpc10*/;
                       Tsp22_SPILL_256 <= 64'sh0;
                       end 
                      
                  13'sd4614/*4614:xpc10*/:  begin 
                       xpc10 <= 13'sd4615/*4615:xpc10*/;
                       Tsco0_2_V_0 <= Tsfl0_9_V_7;
                       end 
                      
                  13'sd4615/*4615:xpc10*/:  begin 
                       xpc10 <= 13'sd4616/*4616:xpc10*/;
                       Tsco0_2_V_1 <= 8'h0;
                       end 
                      
                  13'sd4620/*4620:xpc10*/:  begin 
                       xpc10 <= 13'sd4621/*4621:xpc10*/;
                       Tsco0_2_V_1 <= 8'h20;
                       end 
                      
                  13'sd4624/*4624:xpc10*/:  begin 
                       xpc10 <= 13'sd4625/*4625:xpc10*/;
                       Tsco3_7_V_0 <= rtl_unsigned_bitextract6(64'h_ffff_ffff&Tsco0_2_V_0);
                       end 
                      
                  13'sd4625/*4625:xpc10*/:  begin 
                       xpc10 <= 13'sd4626/*4626:xpc10*/;
                       Tsco3_7_V_1 <= 8'h0;
                       end 
                      
                  13'sd4630/*4630:xpc10*/:  begin 
                       xpc10 <= 13'sd4631/*4631:xpc10*/;
                       Tsco3_7_V_1 <= 8'h10;
                       end 
                      
                  13'sd4631/*4631:xpc10*/:  begin 
                       xpc10 <= 13'sd4632/*4632:xpc10*/;
                       Tsco3_7_V_0 <= (Tsco3_7_V_0<<32'sd16);
                       end 
                      
                  13'sd4639/*4639:xpc10*/:  begin 
                       xpc10 <= 13'sd4640/*4640:xpc10*/;
                       Tsco3_7_V_1 <= rtl_unsigned_bitextract7(8'd8+Tsco3_7_V_1);
                       end 
                      
                  13'sd4640/*4640:xpc10*/:  begin 
                       xpc10 <= 13'sd4641/*4641:xpc10*/;
                       Tsco3_7_V_0 <= (Tsco3_7_V_0<<32'sd8);
                       end 
                      
                  13'sd4644/*4644:xpc10*/:  begin 
                       xpc10 <= 13'sd4645/*4645:xpc10*/;
                       Tsco3_7_V_1 <= rtl_unsigned_bitextract7(Tsco3_7_V_1+A_8_US_CC_SCALbx16_ARA0[$unsigned((Tsco3_7_V_0>>32'sd24))]
                      );

                       end 
                      
                  13'sd4645/*4645:xpc10*/:  begin 
                       xpc10 <= 13'sd4646/*4646:xpc10*/;
                       Tsco0_2_V_1 <= rtl_unsigned_bitextract7(Tsco0_2_V_1+Tsco3_7_V_1);
                       end 
                      
                  13'sd4646/*4646:xpc10*/:  begin 
                       xpc10 <= 13'sd4647/*4647:xpc10*/;
                       Tsno23_4_V_0 <= $unsigned(-32'sd11+rtl_sign_extend8(Tsco0_2_V_1));
                       end 
                      
                  13'sd4647/*4647:xpc10*/:  begin 
                       xpc10 <= 13'sd4648/*4648:xpc10*/;
                       Tsfl0_9_V_7 <= (Tsfl0_9_V_7<<(32'sd63&Tsno23_4_V_0));
                       end 
                      
                  13'sd4648/*4648:xpc10*/:  begin 
                       xpc10 <= 13'sd4649/*4649:xpc10*/;
                       Tsfl0_9_V_4 <= rtl_signed_bitextract0(rtl_sign_extend9(16'sd1)+(0-Tsno23_4_V_0));
                       end 
                      
                  13'sd4652/*4652:xpc10*/:  begin 
                       xpc10 <= 13'sd4653/*4653:xpc10*/;
                       Tsfl0_9_V_5 <= rtl_signed_bitextract0(-16'sd1023+Tsfl0_9_V_3+Tsfl0_9_V_4);
                       end 
                      
                  13'sd4653/*4653:xpc10*/:  begin 
                       xpc10 <= 13'sd4654/*4654:xpc10*/;
                       Tsfl0_9_V_6 <= ((64'sh10_0000_0000_0000|Tsfl0_9_V_6)<<32'sd10);
                       end 
                      
                  13'sd4654/*4654:xpc10*/:  begin 
                       xpc10 <= 13'sd4655/*4655:xpc10*/;
                       Tsfl0_9_V_7 <= ((64'sh10_0000_0000_0000|Tsfl0_9_V_7)<<32'sd11);
                       end 
                      
                  13'sd4655/*4655:xpc10*/:  begin 
                       xpc10 <= 13'sd4656/*4656:xpc10*/;
                       Tsmu24_24_V_1 <= rtl_unsigned_bitextract6(64'h_ffff_ffff&Tsfl0_9_V_6);
                       end 
                      
                  13'sd4656/*4656:xpc10*/:  begin 
                       xpc10 <= 13'sd4657/*4657:xpc10*/;
                       Tsmu24_24_V_0 <= rtl_unsigned_bitextract6((Tsfl0_9_V_6>>32'sd32));
                       end 
                      
                  13'sd4657/*4657:xpc10*/:  begin 
                       xpc10 <= 13'sd4658/*4658:xpc10*/;
                       Tsmu24_24_V_3 <= rtl_unsigned_bitextract6(64'h_ffff_ffff&Tsfl0_9_V_7);
                       end 
                      
                  13'sd4658/*4658:xpc10*/:  begin 
                       xpc10 <= 13'sd4659/*4659:xpc10*/;
                       Tsmu24_24_V_2 <= rtl_unsigned_bitextract6((Tsfl0_9_V_7>>32'sd32));
                       end 
                      
                  13'sd4659/*4659:xpc10*/:  begin 
                       xpc10 <= 13'sd4660/*4660:xpc10*/;
                       Tsmu24_24_V_7 <= rtl_unsigned_extend10(Tsmu24_24_V_1)*rtl_unsigned_extend10(Tsmu24_24_V_3);
                       end 
                      
                  13'sd4660/*4660:xpc10*/:  begin 
                       xpc10 <= 13'sd4661/*4661:xpc10*/;
                       Tsmu24_24_V_5 <= rtl_unsigned_extend10(Tsmu24_24_V_1)*rtl_unsigned_extend10(Tsmu24_24_V_2);
                       end 
                      
                  13'sd4661/*4661:xpc10*/:  begin 
                       xpc10 <= 13'sd4662/*4662:xpc10*/;
                       Tsmu24_24_V_6 <= rtl_unsigned_extend10(Tsmu24_24_V_0)*rtl_unsigned_extend10(Tsmu24_24_V_3);
                       end 
                      
                  13'sd4662/*4662:xpc10*/:  begin 
                       xpc10 <= 13'sd4663/*4663:xpc10*/;
                       Tsmu24_24_V_4 <= rtl_unsigned_extend10(Tsmu24_24_V_0)*rtl_unsigned_extend10(Tsmu24_24_V_2);
                       end 
                      
                  13'sd4663/*4663:xpc10*/:  begin 
                       xpc10 <= 13'sd4664/*4664:xpc10*/;
                       Tsmu24_24_V_5 <= Tsmu24_24_V_5+Tsmu24_24_V_6;
                       end 
                      
                  13'sd4673/*4673:xpc10*/:  begin 
                       xpc10 <= 13'sd4674/*4674:xpc10*/;
                       fastspilldup18 <= Tsmu24_24_V_4;
                       end 
                      
                  13'sd4674/*4674:xpc10*/:  begin 
                       xpc10 <= 13'sd4675/*4675:xpc10*/;
                       Tsm24_SPILL_264 <= fastspilldup18;
                       end 
                      
                  13'sd4675/*4675:xpc10*/:  begin 
                       xpc10 <= 13'sd4676/*4676:xpc10*/;
                       Tsm24_SPILL_257 <= fastspilldup18;
                       end 
                      
                  13'sd4680/*4680:xpc10*/:  begin 
                       xpc10 <= 13'sd4681/*4681:xpc10*/;
                       Tsm24_SPILL_259 <= 64'sh1;
                       end 
                      
                  13'sd4681/*4681:xpc10*/:  begin 
                       xpc10 <= 13'sd4682/*4682:xpc10*/;
                       Tsm24_SPILL_258 <= Tsm24_SPILL_257;
                       end 
                      
                  13'sd4685/*4685:xpc10*/:  begin 
                       xpc10 <= 13'sd4686/*4686:xpc10*/;
                       Tsmu24_24_V_4 <= Tsm24_SPILL_258+(Tsm24_SPILL_259<<32'sd32)+(Tsmu24_24_V_5>>32'sd32);
                       end 
                      
                  13'sd4686/*4686:xpc10*/:  begin 
                       xpc10 <= 13'sd4687/*4687:xpc10*/;
                       Tsmu24_24_V_5 <= (Tsmu24_24_V_5<<32'sd32);
                       end 
                      
                  13'sd4687/*4687:xpc10*/:  begin 
                       xpc10 <= 13'sd4688/*4688:xpc10*/;
                       Tsmu24_24_V_7 <= Tsmu24_24_V_7+Tsmu24_24_V_5;
                       end 
                      
                  13'sd4688/*4688:xpc10*/:  begin 
                       xpc10 <= 13'sd4689/*4689:xpc10*/;
                       fastspilldup20 <= Tsmu24_24_V_4;
                       end 
                      
                  13'sd4689/*4689:xpc10*/:  begin 
                       xpc10 <= 13'sd4690/*4690:xpc10*/;
                       Tsm24_SPILL_263 <= fastspilldup20;
                       end 
                      
                  13'sd4690/*4690:xpc10*/:  begin 
                       xpc10 <= 13'sd4691/*4691:xpc10*/;
                       Tsm24_SPILL_260 <= fastspilldup20;
                       end 
                      
                  13'sd4695/*4695:xpc10*/:  begin 
                       xpc10 <= 13'sd4696/*4696:xpc10*/;
                       Tsm24_SPILL_262 <= 64'sh1;
                       end 
                      
                  13'sd4696/*4696:xpc10*/:  begin 
                       xpc10 <= 13'sd4697/*4697:xpc10*/;
                       Tsm24_SPILL_261 <= Tsm24_SPILL_260;
                       end 
                      
                  13'sd4700/*4700:xpc10*/:  begin 
                       xpc10 <= 13'sd4701/*4701:xpc10*/;
                       Tsmu24_24_V_4 <= Tsm24_SPILL_262+Tsm24_SPILL_261;
                       end 
                      
                  13'sd4701/*4701:xpc10*/:  begin 
                       xpc10 <= 13'sd4702/*4702:xpc10*/;
                       Tsfl0_9_V_9 <= Tsmu24_24_V_7;
                       end 
                      
                  13'sd4702/*4702:xpc10*/:  begin 
                       xpc10 <= 13'sd4703/*4703:xpc10*/;
                       Tsfl0_9_V_8 <= Tsmu24_24_V_4;
                       end 
                      
                  13'sd4703/*4703:xpc10*/:  begin 
                       xpc10 <= 13'sd4704/*4704:xpc10*/;
                       fastspilldup22 <= Tsfl0_9_V_8;
                       end 
                      
                  13'sd4704/*4704:xpc10*/:  begin 
                       xpc10 <= 13'sd4705/*4705:xpc10*/;
                       Tsf0_SPILL_260 <= fastspilldup22;
                       end 
                      
                  13'sd4705/*4705:xpc10*/:  begin 
                       xpc10 <= 13'sd4706/*4706:xpc10*/;
                       Tsf0_SPILL_257 <= fastspilldup22;
                       end 
                      endcase
              if ((Tsfl1_8_V_9==32'sd0/*0:Tsfl1.8_V_9*/))  begin if ((13'sd4137/*4137:xpc10*/==xpc10))  xpc10 <= 13'sd4326/*4326:xpc10*/;
                       end 
                   else if ((13'sd4137/*4137:xpc10*/==xpc10))  xpc10 <= 13'sd4138/*4138:xpc10*/;
                      
              case (xpc10)
                  13'sd3519/*3519:xpc10*/:  begin 
                       xpc10 <= 13'sd3520/*3520:xpc10*/;
                       Tsf1SPILL10_259 <= 64'sh1;
                       end 
                      
                  13'sd3520/*3520:xpc10*/:  begin 
                       xpc10 <= 13'sd3521/*3521:xpc10*/;
                       Tsf1SPILL10_258 <= Tsf1SPILL10_257;
                       end 
                      
                  13'sd3524/*3524:xpc10*/:  begin 
                       xpc10 <= 13'sd3525/*3525:xpc10*/;
                       Tsfl1_24_V_8 <= Tsf1SPILL10_259|Tsf1SPILL10_258;
                       end 
                      
                  13'sd3525/*3525:xpc10*/: if (((Tsfl1_24_V_8<<32'sd1)<64'sh0))  xpc10 <= 13'sd3532/*3532:xpc10*/;
                       else  xpc10 <= 13'sd3526/*3526:xpc10*/;

                  13'sd3529/*3529:xpc10*/:  begin 
                       xpc10 <= 13'sd3530/*3530:xpc10*/;
                       Tsfl1_24_V_8 <= (Tsfl1_24_V_8<<32'sd1);
                       end 
                      
                  13'sd3530/*3530:xpc10*/:  begin 
                       xpc10 <= 13'sd3531/*3531:xpc10*/;
                       Tsfl1_24_V_5 <= rtl_signed_bitextract0(-16'sd1+Tsfl1_24_V_5);
                       end 
                      
                  13'sd3534/*3534:xpc10*/:  begin 
                       xpc10 <= 13'sd3535/*3535:xpc10*/;
                       Tsro29_4_V_0 <= rtl_signed_bitextract0(Tsfl1_24_V_5);
                       end 
                      
                  13'sd3535/*3535:xpc10*/:  begin 
                       xpc10 <= 13'sd3536/*3536:xpc10*/;
                       Tsro29_4_V_1 <= Tsfl1_24_V_8;
                       end 
                      
                  13'sd3538/*3538:xpc10*/:  begin 
                       xpc10 <= 13'sd3539/*3539:xpc10*/;
                       Tsro29_4_V_5 <= 16'sh200;
                       end 
                      
                  13'sd3542/*3542:xpc10*/:  begin 
                       xpc10 <= 13'sd3543/*3543:xpc10*/;
                       Tsro29_4_V_6 <= rtl_signed_bitextract2(64'sh3ff&Tsro29_4_V_1);
                       end 
                      
                  13'sd3564/*3564:xpc10*/:  begin 
                       xpc10 <= 13'sd3565/*3565:xpc10*/;
                       Tsp13_SPILL_256 <= 64'sh1;
                       end 
                      
                  13'sd3568/*3568:xpc10*/:  begin 
                       xpc10 <= 13'sd3569/*3569:xpc10*/;
                       fastspilldup44 <= $signed(64'sh_7ff0_0000_0000_0000+(Tsp13_SPILL_256<<32'sd63));
                       end 
                      
                  13'sd3569/*3569:xpc10*/:  begin 
                       xpc10 <= 13'sd3570/*3570:xpc10*/;
                       Tsr29_SPILL_260 <= fastspilldup44;
                       end 
                      
                  13'sd3570/*3570:xpc10*/:  begin 
                       xpc10 <= 13'sd3571/*3571:xpc10*/;
                       Tsr29_SPILL_256 <= fastspilldup44;
                       end 
                      
                  13'sd3575/*3575:xpc10*/:  begin 
                       xpc10 <= 13'sd3576/*3576:xpc10*/;
                       Tsr29_SPILL_258 <= 64'sh1;
                       end 
                      
                  13'sd3576/*3576:xpc10*/:  begin 
                       xpc10 <= 13'sd3577/*3577:xpc10*/;
                       Tsr29_SPILL_257 <= Tsr29_SPILL_256;
                       end 
                      
                  13'sd3580/*3580:xpc10*/:  begin 
                       xpc10 <= 13'sd3581/*3581:xpc10*/;
                       Tsr29_SPILL_259 <= Tsr29_SPILL_257+(0-Tsr29_SPILL_258);
                       end 
                      
                  13'sd3584/*3584:xpc10*/:  begin 
                       xpc10 <= 13'sd3585/*3585:xpc10*/;
                       Tsf1SPILL10_256 <= Tsr29_SPILL_259;
                       end 
                      
                  13'sd3588/*3588:xpc10*/:  begin 
                       xpc10 <= 13'sd3589/*3589:xpc10*/;
                       Tsr29_SPILL_258 <= 64'sh0;
                       end 
                      
                  13'sd3589/*3589:xpc10*/:  begin 
                       xpc10 <= 13'sd3590/*3590:xpc10*/;
                       Tsr29_SPILL_257 <= Tsr29_SPILL_260;
                       end 
                      
                  13'sd3593/*3593:xpc10*/:  begin 
                       xpc10 <= 13'sd3594/*3594:xpc10*/;
                       Tsp13_SPILL_256 <= 64'sh0;
                       end 
                      
                  13'sd3606/*3606:xpc10*/:  begin 
                       xpc10 <= 13'sd3607/*3607:xpc10*/;
                       Tssh18_7_V_0 <= Tsro29_4_V_1;
                       end 
                      
                  13'sd3610/*3610:xpc10*/:  begin 
                       xpc10 <= 13'sd3611/*3611:xpc10*/;
                       Tsro29_4_V_1 <= Tssh18_7_V_0;
                       end 
                      
                  13'sd3611/*3611:xpc10*/:  begin 
                       xpc10 <= 13'sd3612/*3612:xpc10*/;
                       Tsro29_4_V_0 <= 16'sh0;
                       end 
                      
                  13'sd3612/*3612:xpc10*/:  begin 
                       xpc10 <= 13'sd3613/*3613:xpc10*/;
                       Tsro29_4_V_6 <= rtl_signed_bitextract2(64'sh3ff&Tsro29_4_V_1);
                       end 
                      
                  13'sd3632/*3632:xpc10*/:  begin 
                       xpc10 <= 13'sd3633/*3633:xpc10*/;
                       Tsro29_4_V_1 <= (Tsro29_4_V_1+rtl_sign_extend1(Tsro29_4_V_5)>>32'sd10);
                       end 
                      
                  13'sd3637/*3637:xpc10*/:  begin 
                       xpc10 <= 13'sd3638/*3638:xpc10*/;
                       Tsro29_4_V_1 <= -64'sh2&Tsro29_4_V_1;
                       end 
                      
                  13'sd3645/*3645:xpc10*/:  begin 
                       xpc10 <= 13'sd3646/*3646:xpc10*/;
                       Tsro29_4_V_0 <= 16'sh0;
                       end 
                      
                  13'sd3653/*3653:xpc10*/:  begin 
                       xpc10 <= 13'sd3654/*3654:xpc10*/;
                       Tsp27_SPILL_256 <= 64'sh1;
                       end 
                      
                  13'sd3657/*3657:xpc10*/:  begin 
                       xpc10 <= 13'sd3658/*3658:xpc10*/;
                       Tsr29_SPILL_259 <= Tsro29_4_V_1+(Tsp27_SPILL_256<<32'sd63)+(rtl_sign_extend1(Tsro29_4_V_0)<<32'sd52);
                       end 
                      
                  13'sd3661/*3661:xpc10*/:  begin 
                       xpc10 <= 13'sd3662/*3662:xpc10*/;
                       Tsp27_SPILL_256 <= 64'sh0;
                       end 
                      
                  13'sd3669/*3669:xpc10*/:  begin 
                       xpc10 <= 13'sd3670/*3670:xpc10*/;
                       fastspilldup46 <= (Tsro29_4_V_1>>(32'sd63&rtl_signed_bitextract0((0-Tsro29_4_V_0))));
                       end 
                      
                  13'sd3670/*3670:xpc10*/:  begin 
                       xpc10 <= 13'sd3671/*3671:xpc10*/;
                       Tss18_SPILL_259 <= fastspilldup46;
                       end 
                      
                  13'sd3671/*3671:xpc10*/:  begin 
                       xpc10 <= 13'sd3672/*3672:xpc10*/;
                       Tss18_SPILL_256 <= fastspilldup46;
                       end 
                      
                  13'sd3676/*3676:xpc10*/:  begin 
                       xpc10 <= 13'sd3677/*3677:xpc10*/;
                       Tss18_SPILL_258 <= 64'sh1;
                       end 
                      
                  13'sd3677/*3677:xpc10*/:  begin 
                       xpc10 <= 13'sd3678/*3678:xpc10*/;
                       Tss18_SPILL_257 <= Tss18_SPILL_256;
                       end 
                      
                  13'sd3681/*3681:xpc10*/:  begin 
                       xpc10 <= 13'sd3682/*3682:xpc10*/;
                       Tssh18_7_V_0 <= Tss18_SPILL_258|Tss18_SPILL_257;
                       end 
                      
                  13'sd3685/*3685:xpc10*/:  begin 
                       xpc10 <= 13'sd3686/*3686:xpc10*/;
                       Tss18_SPILL_258 <= 64'sh0;
                       end 
                      
                  13'sd3686/*3686:xpc10*/:  begin 
                       xpc10 <= 13'sd3687/*3687:xpc10*/;
                       Tss18_SPILL_257 <= Tss18_SPILL_259;
                       end 
                      
                  13'sd3694/*3694:xpc10*/:  begin 
                       xpc10 <= 13'sd3695/*3695:xpc10*/;
                       Tss18_SPILL_260 <= 64'sh1;
                       end 
                      
                  13'sd3698/*3698:xpc10*/:  begin 
                       xpc10 <= 13'sd3699/*3699:xpc10*/;
                       Tssh18_7_V_0 <= Tss18_SPILL_260;
                       end 
                      
                  13'sd3702/*3702:xpc10*/:  begin 
                       xpc10 <= 13'sd3703/*3703:xpc10*/;
                       Tss18_SPILL_260 <= 64'sh0;
                       end 
                      
                  13'sd3706/*3706:xpc10*/:  begin 
                       xpc10 <= 13'sd3707/*3707:xpc10*/;
                       Tsf1SPILL10_259 <= 64'sh0;
                       end 
                      
                  13'sd3707/*3707:xpc10*/:  begin 
                       xpc10 <= 13'sd3708/*3708:xpc10*/;
                       Tsf1SPILL10_258 <= Tsf1SPILL10_260;
                       end 
                      
                  13'sd3711/*3711:xpc10*/:  begin 
                       xpc10 <= 13'sd3712/*3712:xpc10*/;
                       Tsm24_SPILL_262 <= 64'sh0;
                       end 
                      
                  13'sd3712/*3712:xpc10*/:  begin 
                       xpc10 <= 13'sd3713/*3713:xpc10*/;
                       Tsm24_SPILL_261 <= Tsm24_SPILL_263;
                       end 
                      
                  13'sd3716/*3716:xpc10*/:  begin 
                       xpc10 <= 13'sd3717/*3717:xpc10*/;
                       Tsm24_SPILL_259 <= 64'sh0;
                       end 
                      
                  13'sd3717/*3717:xpc10*/:  begin 
                       xpc10 <= 13'sd3718/*3718:xpc10*/;
                       Tsm24_SPILL_258 <= Tsm24_SPILL_264;
                       end 
                      
                  13'sd3725/*3725:xpc10*/:  begin 
                       xpc10 <= 13'sd3726/*3726:xpc10*/;
                       Tsco0_2_V_0 <= (Tsco0_2_V_0>>32'sd32);
                       end 
                      
                  13'sd3729/*3729:xpc10*/:  begin 
                       xpc10 <= 13'sd3730/*3730:xpc10*/;
                       Tsco0_2_V_0 <= (Tsco0_2_V_0>>32'sd32);
                       end 
                      
                  13'sd3733/*3733:xpc10*/:  begin 
                       xpc10 <= 13'sd3734/*3734:xpc10*/;
                       Tse0SPILL10_256 <= 32'sd0;
                       end 
                      
                  13'sd3737/*3737:xpc10*/:  begin 
                       xpc10 <= 13'sd3738/*3738:xpc10*/;
                       Tse0_SPILL_256 <= 32'sd0;
                       end 
                      
                  13'sd3741/*3741:xpc10*/:  begin 
                       xpc10 <= 13'sd3742/*3742:xpc10*/;
                       Tsin1_19_V_0 <= (32'sd2*Tdsi1_5_V_2*(32'sd1+32'sd2*Tdsi1_5_V_2)<32'sd0);
                       end 
                      
                  13'sd3746/*3746:xpc10*/:  begin 
                       xpc10 <= 13'sd3747/*3747:xpc10*/;
                       Tsi1_SPILL_257 <= -32'sd2*Tdsi1_5_V_2*(32'sd1+32'sd2*Tdsi1_5_V_2);
                       end 
                      
                  13'sd3750/*3750:xpc10*/:  begin 
                       xpc10 <= 13'sd3751/*3751:xpc10*/;
                       Tsin1_19_V_1 <= Tsi1_SPILL_257;
                       end 
                      
                  13'sd3751/*3751:xpc10*/:  begin 
                       xpc10 <= 13'sd3752/*3752:xpc10*/;
                       Tsco5_4_V_0 <= Tsin1_19_V_1;
                       end 
                      
                  13'sd3752/*3752:xpc10*/:  begin 
                       xpc10 <= 13'sd3753/*3753:xpc10*/;
                       Tsco5_4_V_1 <= 8'h0;
                       end 
                      
                  13'sd3757/*3757:xpc10*/:  begin 
                       xpc10 <= 13'sd3758/*3758:xpc10*/;
                       Tsco5_4_V_1 <= 8'h10;
                       end 
                      
                  13'sd3758/*3758:xpc10*/:  begin 
                       xpc10 <= 13'sd3759/*3759:xpc10*/;
                       Tsco5_4_V_0 <= (Tsco5_4_V_0<<32'sd16);
                       end 
                      
                  13'sd3766/*3766:xpc10*/:  begin 
                       xpc10 <= 13'sd3767/*3767:xpc10*/;
                       Tsco5_4_V_1 <= rtl_unsigned_bitextract7(8'd8+Tsco5_4_V_1);
                       end 
                      
                  13'sd3767/*3767:xpc10*/:  begin 
                       xpc10 <= 13'sd3768/*3768:xpc10*/;
                       Tsco5_4_V_0 <= (Tsco5_4_V_0<<32'sd8);
                       end 
                      
                  13'sd3771/*3771:xpc10*/:  begin 
                       xpc10 <= 13'sd3772/*3772:xpc10*/;
                       Tsco5_4_V_1 <= rtl_unsigned_bitextract7(Tsco5_4_V_1+A_8_US_CC_SCALbx16_ARA0[$unsigned((Tsco5_4_V_0>>32'sd24))]
                      );

                       end 
                      
                  13'sd3772/*3772:xpc10*/:  begin 
                       xpc10 <= 13'sd3773/*3773:xpc10*/;
                       Tsin1_19_V_3 <= $unsigned(32'sd21+rtl_sign_extend8(Tsco5_4_V_1));
                       end 
                      
                  13'sd3773/*3773:xpc10*/:  begin 
                       xpc10 <= 13'sd3774/*3774:xpc10*/;
                       Tsin1_19_V_2 <= rtl_unsigned_extend10(Tsin1_19_V_1);
                       end 
                      
                  13'sd3778/*3778:xpc10*/:  begin 
                       xpc10 <= 13'sd3779/*3779:xpc10*/;
                       Tsp5_SPILL_256 <= 64'sh1;
                       end 
                      
                  13'sd3782/*3782:xpc10*/:  begin 
                       xpc10 <= 13'sd3783/*3783:xpc10*/;
                       Tsi1_SPILL_256 <= (Tsp5_SPILL_256<<32'sd63)+(rtl_sign_extend11(rtl_signed_bitextract0(rtl_sign_extend9(16'sd1074
                      )+(0-Tsin1_19_V_3)))<<32'sd52)+(Tsin1_19_V_2<<(32'sd63&Tsin1_19_V_3));

                       end 
                      
                  13'sd3786/*3786:xpc10*/:  begin 
                       xpc10 <= 13'sd3787/*3787:xpc10*/;
                       Tsp5_SPILL_256 <= 64'sh0;
                       end 
                      
                  13'sd3790/*3790:xpc10*/:  begin 
                       xpc10 <= 13'sd3791/*3791:xpc10*/;
                       Tsi1_SPILL_257 <= 32'sd2*Tdsi1_5_V_2*(32'sd1+32'sd2*Tdsi1_5_V_2);
                       end 
                      
                  13'sd3798/*3798:xpc10*/:  begin 
                       xpc10 <= 13'sd3799/*3799:xpc10*/;
                       Tsp4_SPILL_256 <= Tspr4_3_V_0;
                       end 
                      
                  13'sd3806/*3806:xpc10*/:  begin 
                       xpc10 <= 13'sd3807/*3807:xpc10*/;
                       Tsp4_SPILL_256 <= Tspr4_3_V_1;
                       end 
                      
                  13'sd3810/*3810:xpc10*/:  begin 
                       xpc10 <= 13'sd3811/*3811:xpc10*/;
                       Tsp4_SPILL_256 <= Tspr4_3_V_0;
                       end 
                      
                  13'sd3814/*3814:xpc10*/:  begin 
                       xpc10 <= 13'sd3815/*3815:xpc10*/;
                       Tsf0SPILL12_256 <= 32'sd0;
                       end 
                      
                  13'sd3818/*3818:xpc10*/:  begin 
                       xpc10 <= 13'sd3819/*3819:xpc10*/;
                       Tsf0SPILL10_256 <= 32'sd0;
                       end 
                      
                  13'sd3831/*3831:xpc10*/:  begin 
                       xpc10 <= 13'sd3832/*3832:xpc10*/;
                       Tsf1_SPILL_256 <= 64'h_7fff_ffff_ffff_ffff;
                       end 
                      
                  13'sd3839/*3839:xpc10*/:  begin 
                       xpc10 <= 13'sd3840/*3840:xpc10*/;
                       Tsp8_SPILL_256 <= 64'sh1;
                       end 
                      
                  13'sd3843/*3843:xpc10*/:  begin 
                       xpc10 <= 13'sd3844/*3844:xpc10*/;
                       Tsf1_SPILL_256 <= $signed(64'sh_7ff0_0000_0000_0000+(Tsp8_SPILL_256<<32'sd63));
                       end 
                      
                  13'sd3847/*3847:xpc10*/:  begin 
                       xpc10 <= 13'sd3848/*3848:xpc10*/;
                       Tsp8_SPILL_256 <= 64'sh0;
                       end 
                      
                  13'sd3859/*3859:xpc10*/:  begin 
                       xpc10 <= 13'sd3860/*3860:xpc10*/;
                       Tspr11_2_V_0 <= Tdsi1_5_V_1;
                       end 
                      
                  13'sd3860/*3860:xpc10*/:  begin 
                       xpc10 <= 13'sd3861/*3861:xpc10*/;
                       Tspr11_2_V_1 <= Tdsi1_5_V_3;
                       end 
                      
                  13'sd3865/*3865:xpc10*/:  begin 
                       xpc10 <= 13'sd3866/*3866:xpc10*/;
                       Tsf0SPILL10_256 <= rtl_sign_extend3((32'sd0/*0:USA26*/==(32'sd0/*0:USA24*/==(64'sh7_ffff_ffff_ffff&Tspr11_2_V_0
                      ))));

                       end 
                      
                  13'sd3869/*3869:xpc10*/:  begin 
                       xpc10 <= 13'sd3870/*3870:xpc10*/;
                       Tspr11_2_V_2 <= rtl_unsigned_bitextract4(Tsf0SPILL10_256);
                       end 
                      
                  13'sd3870/*3870:xpc10*/:  begin 
                       xpc10 <= 13'sd3871/*3871:xpc10*/;
                       Tspr11_2_V_3 <= (32'sd0<rtl_sign_extend5(54'sd9007199254740992)+(Tspr11_2_V_1<<32'sd1));
                       end 
                      
                  13'sd3875/*3875:xpc10*/:  begin 
                       xpc10 <= 13'sd3876/*3876:xpc10*/;
                       Tsf0SPILL12_256 <= rtl_sign_extend3((32'sd0/*0:USA32*/==(32'sd0/*0:USA30*/==(64'sh7_ffff_ffff_ffff&Tspr11_2_V_1
                      ))));

                       end 
                      
                  13'sd3879/*3879:xpc10*/:  begin 
                       xpc10 <= 13'sd3880/*3880:xpc10*/;
                       Tspr11_2_V_4 <= rtl_unsigned_bitextract4(Tsf0SPILL12_256);
                       end 
                      
                  13'sd3880/*3880:xpc10*/:  begin 
                       xpc10 <= 13'sd3881/*3881:xpc10*/;
                       Tspr11_2_V_0 <= 64'sh8_0000_0000_0000|Tspr11_2_V_0;
                       end 
                      
                  13'sd3881/*3881:xpc10*/:  begin 
                       xpc10 <= 13'sd3882/*3882:xpc10*/;
                       Tspr11_2_V_1 <= 64'sh8_0000_0000_0000|Tspr11_2_V_1;
                       end 
                      
                  13'sd3894/*3894:xpc10*/:  begin 
                       xpc10 <= 13'sd3895/*3895:xpc10*/;
                       Tsp11_SPILL_256 <= Tspr11_2_V_1;
                       end 
                      
                  13'sd3898/*3898:xpc10*/:  begin 
                       xpc10 <= 13'sd3899/*3899:xpc10*/;
                       Tsf1_SPILL_256 <= Tsp11_SPILL_256;
                       end 
                      
                  13'sd3906/*3906:xpc10*/:  begin 
                       xpc10 <= 13'sd3907/*3907:xpc10*/;
                       Tsp11_SPILL_256 <= Tspr11_2_V_0;
                       end 
                      
                  13'sd3914/*3914:xpc10*/:  begin 
                       xpc10 <= 13'sd3915/*3915:xpc10*/;
                       Tsp11_SPILL_256 <= Tspr11_2_V_1;
                       end 
                      
                  13'sd3918/*3918:xpc10*/:  begin 
                       xpc10 <= 13'sd3919/*3919:xpc10*/;
                       Tsp11_SPILL_256 <= Tspr11_2_V_0;
                       end 
                      
                  13'sd3922/*3922:xpc10*/:  begin 
                       xpc10 <= 13'sd3923/*3923:xpc10*/;
                       Tsf0SPILL12_256 <= 32'sd0;
                       end 
                      
                  13'sd3926/*3926:xpc10*/:  begin 
                       xpc10 <= 13'sd3927/*3927:xpc10*/;
                       Tsf0SPILL10_256 <= 32'sd0;
                       end 
                      
                  13'sd3939/*3939:xpc10*/:  begin 
                       xpc10 <= 13'sd3940/*3940:xpc10*/;
                       Tsf1_SPILL_256 <= 64'h_7fff_ffff_ffff_ffff;
                       end 
                      
                  13'sd3947/*3947:xpc10*/:  begin 
                       xpc10 <= 13'sd3948/*3948:xpc10*/;
                       Tsp15_SPILL_256 <= 64'sh1;
                       end 
                      
                  13'sd3951/*3951:xpc10*/:  begin 
                       xpc10 <= 13'sd3952/*3952:xpc10*/;
                       Tsf1_SPILL_256 <= $signed(64'sh_7ff0_0000_0000_0000+(Tsp15_SPILL_256<<32'sd63));
                       end 
                      
                  13'sd3955/*3955:xpc10*/:  begin 
                       xpc10 <= 13'sd3956/*3956:xpc10*/;
                       Tsp15_SPILL_256 <= 64'sh0;
                       end 
                      
                  13'sd3971/*3971:xpc10*/:  begin 
                       xpc10 <= 13'sd3972/*3972:xpc10*/;
                       Tsp18_SPILL_256 <= 64'sh1;
                       end 
                      
                  13'sd3975/*3975:xpc10*/:  begin 
                       xpc10 <= 13'sd3976/*3976:xpc10*/;
                       Tsf1_SPILL_256 <= $signed(64'sh0+(Tsp18_SPILL_256<<32'sd63));
                       end 
                      
                  13'sd3979/*3979:xpc10*/:  begin 
                       xpc10 <= 13'sd3980/*3980:xpc10*/;
                       Tsp18_SPILL_256 <= 64'sh0;
                       end 
                      
                  13'sd3983/*3983:xpc10*/:  begin 
                       xpc10 <= 13'sd3984/*3984:xpc10*/;
                       Tsco0_2_V_0 <= Tsfl1_8_V_6;
                       end 
                      
                  13'sd3984/*3984:xpc10*/:  begin 
                       xpc10 <= 13'sd3985/*3985:xpc10*/;
                       Tsco0_2_V_1 <= 8'h0;
                       end 
                      
                  13'sd3989/*3989:xpc10*/:  begin 
                       xpc10 <= 13'sd3990/*3990:xpc10*/;
                       Tsco0_2_V_1 <= 8'h20;
                       end 
                      
                  13'sd3993/*3993:xpc10*/:  begin 
                       xpc10 <= 13'sd3994/*3994:xpc10*/;
                       Tsco3_7_V_0 <= rtl_unsigned_bitextract6(64'h_ffff_ffff&Tsco0_2_V_0);
                       end 
                      
                  13'sd3994/*3994:xpc10*/:  begin 
                       xpc10 <= 13'sd3995/*3995:xpc10*/;
                       Tsco3_7_V_1 <= 8'h0;
                       end 
                      
                  13'sd3999/*3999:xpc10*/:  begin 
                       xpc10 <= 13'sd4000/*4000:xpc10*/;
                       Tsco3_7_V_1 <= 8'h10;
                       end 
                      
                  13'sd4000/*4000:xpc10*/:  begin 
                       xpc10 <= 13'sd4001/*4001:xpc10*/;
                       Tsco3_7_V_0 <= (Tsco3_7_V_0<<32'sd16);
                       end 
                      
                  13'sd4008/*4008:xpc10*/:  begin 
                       xpc10 <= 13'sd4009/*4009:xpc10*/;
                       Tsco3_7_V_1 <= rtl_unsigned_bitextract7(8'd8+Tsco3_7_V_1);
                       end 
                      
                  13'sd4009/*4009:xpc10*/:  begin 
                       xpc10 <= 13'sd4010/*4010:xpc10*/;
                       Tsco3_7_V_0 <= (Tsco3_7_V_0<<32'sd8);
                       end 
                      
                  13'sd4013/*4013:xpc10*/:  begin 
                       xpc10 <= 13'sd4014/*4014:xpc10*/;
                       Tsco3_7_V_1 <= rtl_unsigned_bitextract7(Tsco3_7_V_1+A_8_US_CC_SCALbx16_ARA0[$unsigned((Tsco3_7_V_0>>32'sd24))]
                      );

                       end 
                      
                  13'sd4014/*4014:xpc10*/:  begin 
                       xpc10 <= 13'sd4015/*4015:xpc10*/;
                       Tsco0_2_V_1 <= rtl_unsigned_bitextract7(Tsco0_2_V_1+Tsco3_7_V_1);
                       end 
                      
                  13'sd4015/*4015:xpc10*/:  begin 
                       xpc10 <= 13'sd4016/*4016:xpc10*/;
                       Tsno19_4_V_0 <= $unsigned(-32'sd11+rtl_sign_extend8(Tsco0_2_V_1));
                       end 
                      
                  13'sd4016/*4016:xpc10*/:  begin 
                       xpc10 <= 13'sd4017/*4017:xpc10*/;
                       Tsfl1_8_V_6 <= (Tsfl1_8_V_6<<(32'sd63&Tsno19_4_V_0));
                       end 
                      
                  13'sd4017/*4017:xpc10*/:  begin 
                       xpc10 <= 13'sd4018/*4018:xpc10*/;
                       Tsfl1_8_V_3 <= rtl_signed_bitextract0(rtl_sign_extend9(16'sd1)+(0-Tsno19_4_V_0));
                       end 
                      
                  13'sd4033/*4033:xpc10*/:  begin 
                       xpc10 <= 13'sd4034/*4034:xpc10*/;
                       Tsp22_SPILL_256 <= 64'sh1;
                       end 
                      
                  13'sd4037/*4037:xpc10*/:  begin 
                       xpc10 <= 13'sd4038/*4038:xpc10*/;
                       Tsf1_SPILL_256 <= $signed(64'sh0+(Tsp22_SPILL_256<<32'sd63));
                       end 
                      
                  13'sd4041/*4041:xpc10*/:  begin 
                       xpc10 <= 13'sd4042/*4042:xpc10*/;
                       Tsp22_SPILL_256 <= 64'sh0;
                       end 
                      
                  13'sd4045/*4045:xpc10*/:  begin 
                       xpc10 <= 13'sd4046/*4046:xpc10*/;
                       Tsco0_2_V_0 <= Tsfl1_8_V_7;
                       end 
                      
                  13'sd4046/*4046:xpc10*/:  begin 
                       xpc10 <= 13'sd4047/*4047:xpc10*/;
                       Tsco0_2_V_1 <= 8'h0;
                       end 
                      
                  13'sd4051/*4051:xpc10*/:  begin 
                       xpc10 <= 13'sd4052/*4052:xpc10*/;
                       Tsco0_2_V_1 <= 8'h20;
                       end 
                      
                  13'sd4055/*4055:xpc10*/:  begin 
                       xpc10 <= 13'sd4056/*4056:xpc10*/;
                       Tsco3_7_V_0 <= rtl_unsigned_bitextract6(64'h_ffff_ffff&Tsco0_2_V_0);
                       end 
                      
                  13'sd4056/*4056:xpc10*/:  begin 
                       xpc10 <= 13'sd4057/*4057:xpc10*/;
                       Tsco3_7_V_1 <= 8'h0;
                       end 
                      
                  13'sd4061/*4061:xpc10*/:  begin 
                       xpc10 <= 13'sd4062/*4062:xpc10*/;
                       Tsco3_7_V_1 <= 8'h10;
                       end 
                      
                  13'sd4062/*4062:xpc10*/:  begin 
                       xpc10 <= 13'sd4063/*4063:xpc10*/;
                       Tsco3_7_V_0 <= (Tsco3_7_V_0<<32'sd16);
                       end 
                      
                  13'sd4070/*4070:xpc10*/:  begin 
                       xpc10 <= 13'sd4071/*4071:xpc10*/;
                       Tsco3_7_V_1 <= rtl_unsigned_bitextract7(8'd8+Tsco3_7_V_1);
                       end 
                      
                  13'sd4071/*4071:xpc10*/:  begin 
                       xpc10 <= 13'sd4072/*4072:xpc10*/;
                       Tsco3_7_V_0 <= (Tsco3_7_V_0<<32'sd8);
                       end 
                      
                  13'sd4075/*4075:xpc10*/:  begin 
                       xpc10 <= 13'sd4076/*4076:xpc10*/;
                       Tsco3_7_V_1 <= rtl_unsigned_bitextract7(Tsco3_7_V_1+A_8_US_CC_SCALbx16_ARA0[$unsigned((Tsco3_7_V_0>>32'sd24))]
                      );

                       end 
                      
                  13'sd4076/*4076:xpc10*/:  begin 
                       xpc10 <= 13'sd4077/*4077:xpc10*/;
                       Tsco0_2_V_1 <= rtl_unsigned_bitextract7(Tsco0_2_V_1+Tsco3_7_V_1);
                       end 
                      
                  13'sd4077/*4077:xpc10*/:  begin 
                       xpc10 <= 13'sd4078/*4078:xpc10*/;
                       Tsno23_4_V_0 <= $unsigned(-32'sd11+rtl_sign_extend8(Tsco0_2_V_1));
                       end 
                      
                  13'sd4078/*4078:xpc10*/:  begin 
                       xpc10 <= 13'sd4079/*4079:xpc10*/;
                       Tsfl1_8_V_7 <= (Tsfl1_8_V_7<<(32'sd63&Tsno23_4_V_0));
                       end 
                      
                  13'sd4079/*4079:xpc10*/:  begin 
                       xpc10 <= 13'sd4080/*4080:xpc10*/;
                       Tsfl1_8_V_4 <= rtl_signed_bitextract0(rtl_sign_extend9(16'sd1)+(0-Tsno23_4_V_0));
                       end 
                      
                  13'sd4083/*4083:xpc10*/:  begin 
                       xpc10 <= 13'sd4084/*4084:xpc10*/;
                       Tsfl1_8_V_5 <= rtl_signed_bitextract0(-16'sd1023+Tsfl1_8_V_3+Tsfl1_8_V_4);
                       end 
                      
                  13'sd4084/*4084:xpc10*/:  begin 
                       xpc10 <= 13'sd4085/*4085:xpc10*/;
                       Tsfl1_8_V_6 <= ((64'sh10_0000_0000_0000|Tsfl1_8_V_6)<<32'sd10);
                       end 
                      
                  13'sd4085/*4085:xpc10*/:  begin 
                       xpc10 <= 13'sd4086/*4086:xpc10*/;
                       Tsfl1_8_V_7 <= ((64'sh10_0000_0000_0000|Tsfl1_8_V_7)<<32'sd11);
                       end 
                      
                  13'sd4086/*4086:xpc10*/:  begin 
                       xpc10 <= 13'sd4087/*4087:xpc10*/;
                       Tsmu24_24_V_1 <= rtl_unsigned_bitextract6(64'h_ffff_ffff&Tsfl1_8_V_6);
                       end 
                      
                  13'sd4087/*4087:xpc10*/:  begin 
                       xpc10 <= 13'sd4088/*4088:xpc10*/;
                       Tsmu24_24_V_0 <= rtl_unsigned_bitextract6((Tsfl1_8_V_6>>32'sd32));
                       end 
                      
                  13'sd4088/*4088:xpc10*/:  begin 
                       xpc10 <= 13'sd4089/*4089:xpc10*/;
                       Tsmu24_24_V_3 <= rtl_unsigned_bitextract6(64'h_ffff_ffff&Tsfl1_8_V_7);
                       end 
                      
                  13'sd4089/*4089:xpc10*/:  begin 
                       xpc10 <= 13'sd4090/*4090:xpc10*/;
                       Tsmu24_24_V_2 <= rtl_unsigned_bitextract6((Tsfl1_8_V_7>>32'sd32));
                       end 
                      
                  13'sd4090/*4090:xpc10*/:  begin 
                       xpc10 <= 13'sd4091/*4091:xpc10*/;
                       Tsmu24_24_V_7 <= rtl_unsigned_extend10(Tsmu24_24_V_1)*rtl_unsigned_extend10(Tsmu24_24_V_3);
                       end 
                      
                  13'sd4091/*4091:xpc10*/:  begin 
                       xpc10 <= 13'sd4092/*4092:xpc10*/;
                       Tsmu24_24_V_5 <= rtl_unsigned_extend10(Tsmu24_24_V_1)*rtl_unsigned_extend10(Tsmu24_24_V_2);
                       end 
                      
                  13'sd4092/*4092:xpc10*/:  begin 
                       xpc10 <= 13'sd4093/*4093:xpc10*/;
                       Tsmu24_24_V_6 <= rtl_unsigned_extend10(Tsmu24_24_V_0)*rtl_unsigned_extend10(Tsmu24_24_V_3);
                       end 
                      
                  13'sd4093/*4093:xpc10*/:  begin 
                       xpc10 <= 13'sd4094/*4094:xpc10*/;
                       Tsmu24_24_V_4 <= rtl_unsigned_extend10(Tsmu24_24_V_0)*rtl_unsigned_extend10(Tsmu24_24_V_2);
                       end 
                      
                  13'sd4094/*4094:xpc10*/:  begin 
                       xpc10 <= 13'sd4095/*4095:xpc10*/;
                       Tsmu24_24_V_5 <= Tsmu24_24_V_5+Tsmu24_24_V_6;
                       end 
                      
                  13'sd4104/*4104:xpc10*/:  begin 
                       xpc10 <= 13'sd4105/*4105:xpc10*/;
                       fastspilldup28 <= Tsmu24_24_V_4;
                       end 
                      
                  13'sd4105/*4105:xpc10*/:  begin 
                       xpc10 <= 13'sd4106/*4106:xpc10*/;
                       Tsm24_SPILL_264 <= fastspilldup28;
                       end 
                      
                  13'sd4106/*4106:xpc10*/:  begin 
                       xpc10 <= 13'sd4107/*4107:xpc10*/;
                       Tsm24_SPILL_257 <= fastspilldup28;
                       end 
                      
                  13'sd4111/*4111:xpc10*/:  begin 
                       xpc10 <= 13'sd4112/*4112:xpc10*/;
                       Tsm24_SPILL_259 <= 64'sh1;
                       end 
                      
                  13'sd4112/*4112:xpc10*/:  begin 
                       xpc10 <= 13'sd4113/*4113:xpc10*/;
                       Tsm24_SPILL_258 <= Tsm24_SPILL_257;
                       end 
                      
                  13'sd4116/*4116:xpc10*/:  begin 
                       xpc10 <= 13'sd4117/*4117:xpc10*/;
                       Tsmu24_24_V_4 <= Tsm24_SPILL_258+(Tsm24_SPILL_259<<32'sd32)+(Tsmu24_24_V_5>>32'sd32);
                       end 
                      
                  13'sd4117/*4117:xpc10*/:  begin 
                       xpc10 <= 13'sd4118/*4118:xpc10*/;
                       Tsmu24_24_V_5 <= (Tsmu24_24_V_5<<32'sd32);
                       end 
                      
                  13'sd4118/*4118:xpc10*/:  begin 
                       xpc10 <= 13'sd4119/*4119:xpc10*/;
                       Tsmu24_24_V_7 <= Tsmu24_24_V_7+Tsmu24_24_V_5;
                       end 
                      
                  13'sd4119/*4119:xpc10*/:  begin 
                       xpc10 <= 13'sd4120/*4120:xpc10*/;
                       fastspilldup30 <= Tsmu24_24_V_4;
                       end 
                      
                  13'sd4120/*4120:xpc10*/:  begin 
                       xpc10 <= 13'sd4121/*4121:xpc10*/;
                       Tsm24_SPILL_263 <= fastspilldup30;
                       end 
                      
                  13'sd4121/*4121:xpc10*/:  begin 
                       xpc10 <= 13'sd4122/*4122:xpc10*/;
                       Tsm24_SPILL_260 <= fastspilldup30;
                       end 
                      
                  13'sd4126/*4126:xpc10*/:  begin 
                       xpc10 <= 13'sd4127/*4127:xpc10*/;
                       Tsm24_SPILL_262 <= 64'sh1;
                       end 
                      
                  13'sd4127/*4127:xpc10*/:  begin 
                       xpc10 <= 13'sd4128/*4128:xpc10*/;
                       Tsm24_SPILL_261 <= Tsm24_SPILL_260;
                       end 
                      
                  13'sd4131/*4131:xpc10*/:  begin 
                       xpc10 <= 13'sd4132/*4132:xpc10*/;
                       Tsmu24_24_V_4 <= Tsm24_SPILL_262+Tsm24_SPILL_261;
                       end 
                      
                  13'sd4132/*4132:xpc10*/:  begin 
                       xpc10 <= 13'sd4133/*4133:xpc10*/;
                       Tsfl1_8_V_9 <= Tsmu24_24_V_7;
                       end 
                      
                  13'sd4133/*4133:xpc10*/:  begin 
                       xpc10 <= 13'sd4134/*4134:xpc10*/;
                       Tsfl1_8_V_8 <= Tsmu24_24_V_4;
                       end 
                      
                  13'sd4134/*4134:xpc10*/:  begin 
                       xpc10 <= 13'sd4135/*4135:xpc10*/;
                       fastspilldup32 <= Tsfl1_8_V_8;
                       end 
                      
                  13'sd4135/*4135:xpc10*/:  begin 
                       xpc10 <= 13'sd4136/*4136:xpc10*/;
                       Tsf1_SPILL_260 <= fastspilldup32;
                       end 
                      
                  13'sd4136/*4136:xpc10*/:  begin 
                       xpc10 <= 13'sd4137/*4137:xpc10*/;
                       Tsf1_SPILL_257 <= fastspilldup32;
                       end 
                      endcase
              if ((Tsfl1_24_V_9==32'sd0/*0:Tsfl1.24_V_9*/))  begin if ((13'sd3515/*3515:xpc10*/==xpc10))  xpc10 <= 13'sd3704/*3704:xpc10*/;
                       end 
                   else if ((13'sd3515/*3515:xpc10*/==xpc10))  xpc10 <= 13'sd3516/*3516:xpc10*/;
                      
              case (xpc10)
                  13'sd2875/*2875:xpc10*/:  begin 
                       xpc10 <= 13'sd2876/*2876:xpc10*/;
                       Tss18_SPILL_258 <= 64'sh1;
                       end 
                      
                  13'sd2876/*2876:xpc10*/:  begin 
                       xpc10 <= 13'sd2877/*2877:xpc10*/;
                       Tss18_SPILL_257 <= Tss18_SPILL_256;
                       end 
                      
                  13'sd2880/*2880:xpc10*/:  begin 
                       xpc10 <= 13'sd2881/*2881:xpc10*/;
                       Tssh18_7_V_0 <= Tss18_SPILL_258|Tss18_SPILL_257;
                       end 
                      
                  13'sd2884/*2884:xpc10*/:  begin 
                       xpc10 <= 13'sd2885/*2885:xpc10*/;
                       Tss18_SPILL_258 <= 64'sh0;
                       end 
                      
                  13'sd2885/*2885:xpc10*/:  begin 
                       xpc10 <= 13'sd2886/*2886:xpc10*/;
                       Tss18_SPILL_257 <= Tss18_SPILL_259;
                       end 
                      
                  13'sd2893/*2893:xpc10*/:  begin 
                       xpc10 <= 13'sd2894/*2894:xpc10*/;
                       Tss18_SPILL_260 <= 64'sh1;
                       end 
                      
                  13'sd2897/*2897:xpc10*/:  begin 
                       xpc10 <= 13'sd2898/*2898:xpc10*/;
                       Tssh18_7_V_0 <= Tss18_SPILL_260;
                       end 
                      
                  13'sd2901/*2901:xpc10*/:  begin 
                       xpc10 <= 13'sd2902/*2902:xpc10*/;
                       Tss18_SPILL_260 <= 64'sh0;
                       end 
                      
                  13'sd2905/*2905:xpc10*/:  begin 
                       xpc10 <= 13'sd2906/*2906:xpc10*/;
                       Tsf1SPILL12_259 <= 64'sh0;
                       end 
                      
                  13'sd2906/*2906:xpc10*/:  begin 
                       xpc10 <= 13'sd2907/*2907:xpc10*/;
                       Tsf1SPILL12_258 <= Tsf1SPILL12_260;
                       end 
                      
                  13'sd2910/*2910:xpc10*/:  begin 
                       xpc10 <= 13'sd2911/*2911:xpc10*/;
                       Tsfl1_35_V_8 <= -64'd1+Tsfl1_35_V_8;
                       end 
                      
                  13'sd2911/*2911:xpc10*/:  begin 
                       xpc10 <= 13'sd2912/*2912:xpc10*/;
                       Tsad27_13_V_0 <= Tsfl1_35_V_7+Tsfl1_35_V_10;
                       end 
                      
                  13'sd2912/*2912:xpc10*/:  begin 
                       xpc10 <= 13'sd2913/*2913:xpc10*/;
                       Tsfl1_35_V_10 <= Tsad27_13_V_0;
                       end 
                      
                  13'sd2913/*2913:xpc10*/:  begin 
                       xpc10 <= 13'sd2914/*2914:xpc10*/;
                       fastspilldup64 <= 64'sh0+Tsfl1_35_V_9;
                       end 
                      
                  13'sd2914/*2914:xpc10*/:  begin 
                       xpc10 <= 13'sd2915/*2915:xpc10*/;
                       Tsa27_SPILL_262 <= fastspilldup64;
                       end 
                      
                  13'sd2915/*2915:xpc10*/:  begin 
                       xpc10 <= 13'sd2916/*2916:xpc10*/;
                       Tsa27_SPILL_257 <= fastspilldup64;
                       end 
                      
                  13'sd2916/*2916:xpc10*/: if ((Tsad27_13_V_0<Tsfl1_35_V_10))  xpc10 <= 13'sd2917/*2917:xpc10*/;
                       else  xpc10 <= 13'sd2927/*2927:xpc10*/;

                  13'sd2920/*2920:xpc10*/:  begin 
                       xpc10 <= 13'sd2921/*2921:xpc10*/;
                       Tsa27_SPILL_260 <= 64'sh1;
                       end 
                      
                  13'sd2921/*2921:xpc10*/:  begin 
                       xpc10 <= 13'sd2922/*2922:xpc10*/;
                       Tsa27_SPILL_259 <= Tsa27_SPILL_257;
                       end 
                      
                  13'sd2925/*2925:xpc10*/:  begin 
                       xpc10 <= 13'sd2926/*2926:xpc10*/;
                       Tsfl1_35_V_9 <= Tsa27_SPILL_260+Tsa27_SPILL_259;
                       end 
                      
                  13'sd2929/*2929:xpc10*/:  begin 
                       xpc10 <= 13'sd2930/*2930:xpc10*/;
                       Tsa27_SPILL_260 <= 64'sh0;
                       end 
                      
                  13'sd2930/*2930:xpc10*/:  begin 
                       xpc10 <= 13'sd2931/*2931:xpc10*/;
                       Tsa27_SPILL_259 <= Tsa27_SPILL_262;
                       end 
                      
                  13'sd2934/*2934:xpc10*/:  begin 
                       xpc10 <= 13'sd2935/*2935:xpc10*/;
                       Tss26_SPILL_260 <= 64'sh0;
                       end 
                      
                  13'sd2935/*2935:xpc10*/:  begin 
                       xpc10 <= 13'sd2936/*2936:xpc10*/;
                       Tss26_SPILL_259 <= Tss26_SPILL_262;
                       end 
                      
                  13'sd2939/*2939:xpc10*/:  begin 
                       xpc10 <= 13'sd2940/*2940:xpc10*/;
                       Tsm26_SPILL_262 <= 64'sh0;
                       end 
                      
                  13'sd2940/*2940:xpc10*/:  begin 
                       xpc10 <= 13'sd2941/*2941:xpc10*/;
                       Tsm26_SPILL_261 <= Tsm26_SPILL_263;
                       end 
                      
                  13'sd2944/*2944:xpc10*/:  begin 
                       xpc10 <= 13'sd2945/*2945:xpc10*/;
                       Tsm26_SPILL_259 <= 64'sh0;
                       end 
                      
                  13'sd2945/*2945:xpc10*/:  begin 
                       xpc10 <= 13'sd2946/*2946:xpc10*/;
                       Tsm26_SPILL_258 <= Tsm26_SPILL_264;
                       end 
                      
                  13'sd2953/*2953:xpc10*/:  begin 
                       xpc10 <= 13'sd2954/*2954:xpc10*/;
                       Tses25_5_V_0 <= (Tsfl1_35_V_7>>32'sd32);
                       end 
                      
                  13'sd2954/*2954:xpc10*/: if ((Tsfl1_35_V_6<(Tses25_5_V_0<<32'sd32)))  xpc10 <= 13'sd3097/*3097:xpc10*/;
                       else  xpc10 <= 13'sd2955/*2955:xpc10*/;

                  13'sd2958/*2958:xpc10*/:  begin 
                       xpc10 <= 13'sd2959/*2959:xpc10*/;
                       Tse25_SPILL_257 <= 64'h_ffff_ffff_0000_0000;
                       end 
                      
                  13'sd2962/*2962:xpc10*/:  begin 
                       xpc10 <= 13'sd2963/*2963:xpc10*/;
                       Tses25_5_V_6 <= Tse25_SPILL_257;
                       end 
                      
                  13'sd2963/*2963:xpc10*/:  begin 
                       xpc10 <= 13'sd2964/*2964:xpc10*/;
                       Tsmu5_7_V_1 <= rtl_unsigned_bitextract6(64'h_ffff_ffff&Tsfl1_35_V_7);
                       end 
                      
                  13'sd2964/*2964:xpc10*/:  begin 
                       xpc10 <= 13'sd2965/*2965:xpc10*/;
                       Tsmu5_7_V_0 <= rtl_unsigned_bitextract6((Tsfl1_35_V_7>>32'sd32));
                       end 
                      
                  13'sd2965/*2965:xpc10*/:  begin 
                       xpc10 <= 13'sd2966/*2966:xpc10*/;
                       Tsmu5_7_V_3 <= rtl_unsigned_bitextract6(64'h_ffff_ffff&Tses25_5_V_6);
                       end 
                      
                  13'sd2966/*2966:xpc10*/:  begin 
                       xpc10 <= 13'sd2967/*2967:xpc10*/;
                       Tsmu5_7_V_2 <= rtl_unsigned_bitextract6((Tses25_5_V_6>>32'sd32));
                       end 
                      
                  13'sd2967/*2967:xpc10*/:  begin 
                       xpc10 <= 13'sd2968/*2968:xpc10*/;
                       Tsmu5_7_V_7 <= rtl_unsigned_extend10(Tsmu5_7_V_1)*rtl_unsigned_extend10(Tsmu5_7_V_3);
                       end 
                      
                  13'sd2968/*2968:xpc10*/:  begin 
                       xpc10 <= 13'sd2969/*2969:xpc10*/;
                       Tsmu5_7_V_5 <= rtl_unsigned_extend10(Tsmu5_7_V_1)*rtl_unsigned_extend10(Tsmu5_7_V_2);
                       end 
                      
                  13'sd2969/*2969:xpc10*/:  begin 
                       xpc10 <= 13'sd2970/*2970:xpc10*/;
                       Tsmu5_7_V_6 <= rtl_unsigned_extend10(Tsmu5_7_V_0)*rtl_unsigned_extend10(Tsmu5_7_V_3);
                       end 
                      
                  13'sd2970/*2970:xpc10*/:  begin 
                       xpc10 <= 13'sd2971/*2971:xpc10*/;
                       Tsmu5_7_V_4 <= rtl_unsigned_extend10(Tsmu5_7_V_0)*rtl_unsigned_extend10(Tsmu5_7_V_2);
                       end 
                      
                  13'sd2971/*2971:xpc10*/:  begin 
                       xpc10 <= 13'sd2972/*2972:xpc10*/;
                       Tsmu5_7_V_5 <= Tsmu5_7_V_5+Tsmu5_7_V_6;
                       end 
                      
                  13'sd2981/*2981:xpc10*/:  begin 
                       xpc10 <= 13'sd2982/*2982:xpc10*/;
                       fastspilldup48 <= Tsmu5_7_V_4;
                       end 
                      
                  13'sd2982/*2982:xpc10*/:  begin 
                       xpc10 <= 13'sd2983/*2983:xpc10*/;
                       Tsm5_SPILL_264 <= fastspilldup48;
                       end 
                      
                  13'sd2983/*2983:xpc10*/:  begin 
                       xpc10 <= 13'sd2984/*2984:xpc10*/;
                       Tsm5_SPILL_257 <= fastspilldup48;
                       end 
                      
                  13'sd2988/*2988:xpc10*/:  begin 
                       xpc10 <= 13'sd2989/*2989:xpc10*/;
                       Tsm5_SPILL_259 <= 64'sh1;
                       end 
                      
                  13'sd2989/*2989:xpc10*/:  begin 
                       xpc10 <= 13'sd2990/*2990:xpc10*/;
                       Tsm5_SPILL_258 <= Tsm5_SPILL_257;
                       end 
                      
                  13'sd2993/*2993:xpc10*/:  begin 
                       xpc10 <= 13'sd2994/*2994:xpc10*/;
                       Tsmu5_7_V_4 <= Tsm5_SPILL_258+(Tsm5_SPILL_259<<32'sd32)+(Tsmu5_7_V_5>>32'sd32);
                       end 
                      
                  13'sd2994/*2994:xpc10*/:  begin 
                       xpc10 <= 13'sd2995/*2995:xpc10*/;
                       Tsmu5_7_V_5 <= (Tsmu5_7_V_5<<32'sd32);
                       end 
                      
                  13'sd2995/*2995:xpc10*/:  begin 
                       xpc10 <= 13'sd2996/*2996:xpc10*/;
                       Tsmu5_7_V_7 <= Tsmu5_7_V_7+Tsmu5_7_V_5;
                       end 
                      
                  13'sd2996/*2996:xpc10*/:  begin 
                       xpc10 <= 13'sd2997/*2997:xpc10*/;
                       fastspilldup50 <= Tsmu5_7_V_4;
                       end 
                      
                  13'sd2997/*2997:xpc10*/:  begin 
                       xpc10 <= 13'sd2998/*2998:xpc10*/;
                       Tsm5_SPILL_263 <= fastspilldup50;
                       end 
                      
                  13'sd2998/*2998:xpc10*/:  begin 
                       xpc10 <= 13'sd2999/*2999:xpc10*/;
                       Tsm5_SPILL_260 <= fastspilldup50;
                       end 
                      
                  13'sd2999/*2999:xpc10*/: if ((Tsmu5_7_V_7<Tsmu5_7_V_5))  xpc10 <= 13'sd3000/*3000:xpc10*/;
                       else  xpc10 <= 13'sd3083/*3083:xpc10*/;

                  13'sd3003/*3003:xpc10*/:  begin 
                       xpc10 <= 13'sd3004/*3004:xpc10*/;
                       Tsm5_SPILL_262 <= 64'sh1;
                       end 
                      
                  13'sd3004/*3004:xpc10*/:  begin 
                       xpc10 <= 13'sd3005/*3005:xpc10*/;
                       Tsm5_SPILL_261 <= Tsm5_SPILL_260;
                       end 
                      
                  13'sd3008/*3008:xpc10*/:  begin 
                       xpc10 <= 13'sd3009/*3009:xpc10*/;
                       Tsmu5_7_V_4 <= Tsm5_SPILL_262+Tsm5_SPILL_261;
                       end 
                      
                  13'sd3009/*3009:xpc10*/:  begin 
                       xpc10 <= 13'sd3010/*3010:xpc10*/;
                       Tses25_5_V_5 <= Tsmu5_7_V_7;
                       end 
                      
                  13'sd3010/*3010:xpc10*/:  begin 
                       xpc10 <= 13'sd3011/*3011:xpc10*/;
                       Tses25_5_V_4 <= Tsmu5_7_V_4;
                       end 
                      
                  13'sd3011/*3011:xpc10*/:  begin 
                       xpc10 <= 13'sd3012/*3012:xpc10*/;
                       Tses25_5_V_3 <= 64'sh0+(0-Tses25_5_V_5);
                       end 
                      
                  13'sd3012/*3012:xpc10*/:  begin 
                       xpc10 <= 13'sd3013/*3013:xpc10*/;
                       fastspilldup52 <= Tsfl1_35_V_6+(0-Tses25_5_V_4);
                       end 
                      
                  13'sd3013/*3013:xpc10*/:  begin 
                       xpc10 <= 13'sd3014/*3014:xpc10*/;
                       Tss5_SPILL_262 <= fastspilldup52;
                       end 
                      
                  13'sd3014/*3014:xpc10*/:  begin 
                       xpc10 <= 13'sd3015/*3015:xpc10*/;
                       Tss5_SPILL_257 <= fastspilldup52;
                       end 
                      
                  13'sd3015/*3015:xpc10*/: if ((64'sh0<Tses25_5_V_5))  xpc10 <= 13'sd3016/*3016:xpc10*/;
                       else  xpc10 <= 13'sd3078/*3078:xpc10*/;

                  13'sd3019/*3019:xpc10*/:  begin 
                       xpc10 <= 13'sd3020/*3020:xpc10*/;
                       Tss5_SPILL_260 <= 64'sh1;
                       end 
                      
                  13'sd3020/*3020:xpc10*/:  begin 
                       xpc10 <= 13'sd3021/*3021:xpc10*/;
                       Tss5_SPILL_259 <= Tss5_SPILL_257;
                       end 
                      
                  13'sd3024/*3024:xpc10*/:  begin 
                       xpc10 <= 13'sd3025/*3025:xpc10*/;
                       Tses25_5_V_2 <= Tss5_SPILL_259+(0-Tss5_SPILL_260);
                       end 
                      
                  13'sd3028/*3028:xpc10*/: if ((Tses25_5_V_2<64'sh0))  xpc10 <= 13'sd3053/*3053:xpc10*/;
                       else  xpc10 <= 13'sd3029/*3029:xpc10*/;

                  13'sd3032/*3032:xpc10*/:  begin 
                       xpc10 <= 13'sd3033/*3033:xpc10*/;
                       Tses25_5_V_2 <= (Tses25_5_V_2<<32'sd32)|(Tses25_5_V_3>>32'sd32);
                       end 
                      
                  13'sd3033/*3033:xpc10*/:  begin 
                       xpc10 <= 13'sd3034/*3034:xpc10*/;
                       fastspilldup56 <= Tses25_5_V_6;
                       end 
                      
                  13'sd3034/*3034:xpc10*/:  begin 
                       xpc10 <= 13'sd3035/*3035:xpc10*/;
                       Tse25_SPILL_261 <= fastspilldup56;
                       end 
                      
                  13'sd3035/*3035:xpc10*/:  begin 
                       xpc10 <= 13'sd3036/*3036:xpc10*/;
                       Tse25_SPILL_258 <= fastspilldup56;
                       end 
                      
                  13'sd3036/*3036:xpc10*/: if ((Tses25_5_V_2<(Tses25_5_V_0<<32'sd32)))  xpc10 <= 13'sd3048/*3048:xpc10*/;
                       else  xpc10 <= 13'sd3037/*3037:xpc10*/;

                  13'sd3040/*3040:xpc10*/:  begin 
                       xpc10 <= 13'sd3041/*3041:xpc10*/;
                       Tse25_SPILL_260 <= 64'h_ffff_ffff;
                       end 
                      
                  13'sd3041/*3041:xpc10*/:  begin 
                       xpc10 <= 13'sd3042/*3042:xpc10*/;
                       Tse25_SPILL_259 <= Tse25_SPILL_258;
                       end 
                      
                  13'sd3045/*3045:xpc10*/:  begin 
                       xpc10 <= 13'sd3046/*3046:xpc10*/;
                       Tses25_5_V_6 <= Tse25_SPILL_260|Tse25_SPILL_259;
                       end 
                      
                  13'sd3046/*3046:xpc10*/:  begin 
                       xpc10 <= 13'sd3047/*3047:xpc10*/;
                       Tse25_SPILL_256 <= Tses25_5_V_6;
                       end 
                      
                  13'sd3050/*3050:xpc10*/:  begin 
                       xpc10 <= 13'sd3051/*3051:xpc10*/;
                       Tse25_SPILL_260 <= (Tses25_5_V_2/Tses25_5_V_0);
                       end 
                      
                  13'sd3051/*3051:xpc10*/:  begin 
                       xpc10 <= 13'sd3052/*3052:xpc10*/;
                       Tse25_SPILL_259 <= Tse25_SPILL_261;
                       end 
                      
                  13'sd3055/*3055:xpc10*/:  begin 
                       xpc10 <= 13'sd3056/*3056:xpc10*/;
                       Tses25_5_V_6 <= -64'sh1_0000_0000+Tses25_5_V_6;
                       end 
                      
                  13'sd3056/*3056:xpc10*/:  begin 
                       xpc10 <= 13'sd3057/*3057:xpc10*/;
                       Tses25_5_V_1 <= (Tsfl1_35_V_7<<32'sd32);
                       end 
                      
                  13'sd3057/*3057:xpc10*/:  begin 
                       xpc10 <= 13'sd3058/*3058:xpc10*/;
                       Tsad6_15_V_0 <= Tses25_5_V_3+Tses25_5_V_1;
                       end 
                      
                  13'sd3058/*3058:xpc10*/:  begin 
                       xpc10 <= 13'sd3059/*3059:xpc10*/;
                       Tses25_5_V_3 <= Tsad6_15_V_0;
                       end 
                      
                  13'sd3059/*3059:xpc10*/:  begin 
                       xpc10 <= 13'sd3060/*3060:xpc10*/;
                       fastspilldup54 <= Tses25_5_V_0+Tses25_5_V_2;
                       end 
                      
                  13'sd3060/*3060:xpc10*/:  begin 
                       xpc10 <= 13'sd3061/*3061:xpc10*/;
                       Tsa6_SPILL_262 <= fastspilldup54;
                       end 
                      
                  13'sd3061/*3061:xpc10*/:  begin 
                       xpc10 <= 13'sd3062/*3062:xpc10*/;
                       Tsa6_SPILL_257 <= fastspilldup54;
                       end 
                      
                  13'sd3062/*3062:xpc10*/: if ((Tsad6_15_V_0<Tses25_5_V_3))  xpc10 <= 13'sd3063/*3063:xpc10*/;
                       else  xpc10 <= 13'sd3073/*3073:xpc10*/;

                  13'sd3066/*3066:xpc10*/:  begin 
                       xpc10 <= 13'sd3067/*3067:xpc10*/;
                       Tsa6_SPILL_260 <= 64'sh1;
                       end 
                      
                  13'sd3067/*3067:xpc10*/:  begin 
                       xpc10 <= 13'sd3068/*3068:xpc10*/;
                       Tsa6_SPILL_259 <= Tsa6_SPILL_257;
                       end 
                      
                  13'sd3071/*3071:xpc10*/:  begin 
                       xpc10 <= 13'sd3072/*3072:xpc10*/;
                       Tses25_5_V_2 <= Tsa6_SPILL_260+Tsa6_SPILL_259;
                       end 
                      
                  13'sd3075/*3075:xpc10*/:  begin 
                       xpc10 <= 13'sd3076/*3076:xpc10*/;
                       Tsa6_SPILL_260 <= 64'sh0;
                       end 
                      
                  13'sd3076/*3076:xpc10*/:  begin 
                       xpc10 <= 13'sd3077/*3077:xpc10*/;
                       Tsa6_SPILL_259 <= Tsa6_SPILL_262;
                       end 
                      
                  13'sd3080/*3080:xpc10*/:  begin 
                       xpc10 <= 13'sd3081/*3081:xpc10*/;
                       Tss5_SPILL_260 <= 64'sh0;
                       end 
                      
                  13'sd3081/*3081:xpc10*/:  begin 
                       xpc10 <= 13'sd3082/*3082:xpc10*/;
                       Tss5_SPILL_259 <= Tss5_SPILL_262;
                       end 
                      
                  13'sd3085/*3085:xpc10*/:  begin 
                       xpc10 <= 13'sd3086/*3086:xpc10*/;
                       Tsm5_SPILL_262 <= 64'sh0;
                       end 
                      
                  13'sd3086/*3086:xpc10*/:  begin 
                       xpc10 <= 13'sd3087/*3087:xpc10*/;
                       Tsm5_SPILL_261 <= Tsm5_SPILL_263;
                       end 
                      
                  13'sd3090/*3090:xpc10*/:  begin 
                       xpc10 <= 13'sd3091/*3091:xpc10*/;
                       Tsm5_SPILL_259 <= 64'sh0;
                       end 
                      
                  13'sd3091/*3091:xpc10*/:  begin 
                       xpc10 <= 13'sd3092/*3092:xpc10*/;
                       Tsm5_SPILL_258 <= Tsm5_SPILL_264;
                       end 
                      
                  13'sd3099/*3099:xpc10*/:  begin 
                       xpc10 <= 13'sd3100/*3100:xpc10*/;
                       Tse25_SPILL_257 <= ((Tsfl1_35_V_6/Tses25_5_V_0)<<32'sd32);
                       end 
                      
                  13'sd3103/*3103:xpc10*/:  begin 
                       xpc10 <= 13'sd3104/*3104:xpc10*/;
                       Tsco0_2_V_0 <= (Tsco0_2_V_0>>32'sd32);
                       end 
                      
                  13'sd3107/*3107:xpc10*/:  begin 
                       xpc10 <= 13'sd3108/*3108:xpc10*/;
                       Tsco0_2_V_0 <= (Tsco0_2_V_0>>32'sd32);
                       end 
                      
                  13'sd3111/*3111:xpc10*/:  begin 
                       xpc10 <= 13'sd3112/*3112:xpc10*/;
                       Tse0SPILL14_256 <= 32'sd0;
                       end 
                      
                  13'sd3115/*3115:xpc10*/:  begin 
                       xpc10 <= 13'sd3116/*3116:xpc10*/;
                       Tse0SPILL12_256 <= 32'sd0;
                       end 
                      
                  13'sd3119/*3119:xpc10*/:  begin 
                       xpc10 <= 13'sd3120/*3120:xpc10*/;
                       Tsin1_34_V_0 <= (32'sd2*Tdsi1_5_V_2*(32'sd1+32'sd2*Tdsi1_5_V_2)<32'sd0);
                       end 
                      
                  13'sd3124/*3124:xpc10*/:  begin 
                       xpc10 <= 13'sd3125/*3125:xpc10*/;
                       Tsi1SPILL10_257 <= -32'sd2*Tdsi1_5_V_2*(32'sd1+32'sd2*Tdsi1_5_V_2);
                       end 
                      
                  13'sd3128/*3128:xpc10*/:  begin 
                       xpc10 <= 13'sd3129/*3129:xpc10*/;
                       Tsin1_34_V_1 <= Tsi1SPILL10_257;
                       end 
                      
                  13'sd3129/*3129:xpc10*/:  begin 
                       xpc10 <= 13'sd3130/*3130:xpc10*/;
                       Tsco5_4_V_0 <= Tsin1_34_V_1;
                       end 
                      
                  13'sd3130/*3130:xpc10*/:  begin 
                       xpc10 <= 13'sd3131/*3131:xpc10*/;
                       Tsco5_4_V_1 <= 8'h0;
                       end 
                      
                  13'sd3135/*3135:xpc10*/:  begin 
                       xpc10 <= 13'sd3136/*3136:xpc10*/;
                       Tsco5_4_V_1 <= 8'h10;
                       end 
                      
                  13'sd3136/*3136:xpc10*/:  begin 
                       xpc10 <= 13'sd3137/*3137:xpc10*/;
                       Tsco5_4_V_0 <= (Tsco5_4_V_0<<32'sd16);
                       end 
                      
                  13'sd3144/*3144:xpc10*/:  begin 
                       xpc10 <= 13'sd3145/*3145:xpc10*/;
                       Tsco5_4_V_1 <= rtl_unsigned_bitextract7(8'd8+Tsco5_4_V_1);
                       end 
                      
                  13'sd3145/*3145:xpc10*/:  begin 
                       xpc10 <= 13'sd3146/*3146:xpc10*/;
                       Tsco5_4_V_0 <= (Tsco5_4_V_0<<32'sd8);
                       end 
                      
                  13'sd3149/*3149:xpc10*/:  begin 
                       xpc10 <= 13'sd3150/*3150:xpc10*/;
                       Tsco5_4_V_1 <= rtl_unsigned_bitextract7(Tsco5_4_V_1+A_8_US_CC_SCALbx16_ARA0[$unsigned((Tsco5_4_V_0>>32'sd24))]
                      );

                       end 
                      
                  13'sd3150/*3150:xpc10*/:  begin 
                       xpc10 <= 13'sd3151/*3151:xpc10*/;
                       Tsin1_34_V_3 <= $unsigned(32'sd21+rtl_sign_extend8(Tsco5_4_V_1));
                       end 
                      
                  13'sd3151/*3151:xpc10*/:  begin 
                       xpc10 <= 13'sd3152/*3152:xpc10*/;
                       Tsin1_34_V_2 <= rtl_unsigned_extend10(Tsin1_34_V_1);
                       end 
                      
                  13'sd3156/*3156:xpc10*/:  begin 
                       xpc10 <= 13'sd3157/*3157:xpc10*/;
                       Tsp5_SPILL_256 <= 64'sh1;
                       end 
                      
                  13'sd3160/*3160:xpc10*/:  begin 
                       xpc10 <= 13'sd3161/*3161:xpc10*/;
                       Tsi1SPILL10_256 <= (Tsp5_SPILL_256<<32'sd63)+(rtl_sign_extend11(rtl_signed_bitextract0(rtl_sign_extend9(16'sd1074
                      )+(0-Tsin1_34_V_3)))<<32'sd52)+(Tsin1_34_V_2<<(32'sd63&Tsin1_34_V_3));

                       end 
                      
                  13'sd3164/*3164:xpc10*/:  begin 
                       xpc10 <= 13'sd3165/*3165:xpc10*/;
                       Tsp5_SPILL_256 <= 64'sh0;
                       end 
                      
                  13'sd3168/*3168:xpc10*/:  begin 
                       xpc10 <= 13'sd3169/*3169:xpc10*/;
                       Tsi1SPILL10_257 <= 32'sd2*Tdsi1_5_V_2*(32'sd1+32'sd2*Tdsi1_5_V_2);
                       end 
                      
                  13'sd3176/*3176:xpc10*/:  begin 
                       xpc10 <= 13'sd3177/*3177:xpc10*/;
                       Tsp4_SPILL_256 <= Tspr4_3_V_0;
                       end 
                      
                  13'sd3184/*3184:xpc10*/:  begin 
                       xpc10 <= 13'sd3185/*3185:xpc10*/;
                       Tsp4_SPILL_256 <= Tspr4_3_V_1;
                       end 
                      
                  13'sd3188/*3188:xpc10*/:  begin 
                       xpc10 <= 13'sd3189/*3189:xpc10*/;
                       Tsp4_SPILL_256 <= Tspr4_3_V_0;
                       end 
                      
                  13'sd3192/*3192:xpc10*/:  begin 
                       xpc10 <= 13'sd3193/*3193:xpc10*/;
                       Tsf0SPILL12_256 <= 32'sd0;
                       end 
                      
                  13'sd3196/*3196:xpc10*/:  begin 
                       xpc10 <= 13'sd3197/*3197:xpc10*/;
                       Tsf0SPILL10_256 <= 32'sd0;
                       end 
                      
                  13'sd3209/*3209:xpc10*/:  begin 
                       xpc10 <= 13'sd3210/*3210:xpc10*/;
                       Tsf1SPILL10_256 <= 64'h_7fff_ffff_ffff_ffff;
                       end 
                      
                  13'sd3217/*3217:xpc10*/:  begin 
                       xpc10 <= 13'sd3218/*3218:xpc10*/;
                       Tsp8_SPILL_256 <= 64'sh1;
                       end 
                      
                  13'sd3221/*3221:xpc10*/:  begin 
                       xpc10 <= 13'sd3222/*3222:xpc10*/;
                       Tsf1SPILL10_256 <= $signed(64'sh_7ff0_0000_0000_0000+(Tsp8_SPILL_256<<32'sd63));
                       end 
                      
                  13'sd3225/*3225:xpc10*/:  begin 
                       xpc10 <= 13'sd3226/*3226:xpc10*/;
                       Tsp8_SPILL_256 <= 64'sh0;
                       end 
                      
                  13'sd3237/*3237:xpc10*/:  begin 
                       xpc10 <= 13'sd3238/*3238:xpc10*/;
                       Tspr11_2_V_0 <= Tdsi1_5_V_1;
                       end 
                      
                  13'sd3238/*3238:xpc10*/:  begin 
                       xpc10 <= 13'sd3239/*3239:xpc10*/;
                       Tspr11_2_V_1 <= Tdsi1_5_V_3;
                       end 
                      
                  13'sd3243/*3243:xpc10*/:  begin 
                       xpc10 <= 13'sd3244/*3244:xpc10*/;
                       Tsf0SPILL10_256 <= rtl_sign_extend3((32'sd0/*0:USA26*/==(32'sd0/*0:USA24*/==(64'sh7_ffff_ffff_ffff&Tspr11_2_V_0
                      ))));

                       end 
                      
                  13'sd3247/*3247:xpc10*/:  begin 
                       xpc10 <= 13'sd3248/*3248:xpc10*/;
                       Tspr11_2_V_2 <= rtl_unsigned_bitextract4(Tsf0SPILL10_256);
                       end 
                      
                  13'sd3248/*3248:xpc10*/:  begin 
                       xpc10 <= 13'sd3249/*3249:xpc10*/;
                       Tspr11_2_V_3 <= (32'sd0<rtl_sign_extend5(54'sd9007199254740992)+(Tspr11_2_V_1<<32'sd1));
                       end 
                      
                  13'sd3253/*3253:xpc10*/:  begin 
                       xpc10 <= 13'sd3254/*3254:xpc10*/;
                       Tsf0SPILL12_256 <= rtl_sign_extend3((32'sd0/*0:USA32*/==(32'sd0/*0:USA30*/==(64'sh7_ffff_ffff_ffff&Tspr11_2_V_1
                      ))));

                       end 
                      
                  13'sd3257/*3257:xpc10*/:  begin 
                       xpc10 <= 13'sd3258/*3258:xpc10*/;
                       Tspr11_2_V_4 <= rtl_unsigned_bitextract4(Tsf0SPILL12_256);
                       end 
                      
                  13'sd3258/*3258:xpc10*/:  begin 
                       xpc10 <= 13'sd3259/*3259:xpc10*/;
                       Tspr11_2_V_0 <= 64'sh8_0000_0000_0000|Tspr11_2_V_0;
                       end 
                      
                  13'sd3259/*3259:xpc10*/:  begin 
                       xpc10 <= 13'sd3260/*3260:xpc10*/;
                       Tspr11_2_V_1 <= 64'sh8_0000_0000_0000|Tspr11_2_V_1;
                       end 
                      
                  13'sd3272/*3272:xpc10*/:  begin 
                       xpc10 <= 13'sd3273/*3273:xpc10*/;
                       Tsp11_SPILL_256 <= Tspr11_2_V_1;
                       end 
                      
                  13'sd3276/*3276:xpc10*/:  begin 
                       xpc10 <= 13'sd3277/*3277:xpc10*/;
                       Tsf1SPILL10_256 <= Tsp11_SPILL_256;
                       end 
                      
                  13'sd3284/*3284:xpc10*/:  begin 
                       xpc10 <= 13'sd3285/*3285:xpc10*/;
                       Tsp11_SPILL_256 <= Tspr11_2_V_0;
                       end 
                      
                  13'sd3292/*3292:xpc10*/:  begin 
                       xpc10 <= 13'sd3293/*3293:xpc10*/;
                       Tsp11_SPILL_256 <= Tspr11_2_V_1;
                       end 
                      
                  13'sd3296/*3296:xpc10*/:  begin 
                       xpc10 <= 13'sd3297/*3297:xpc10*/;
                       Tsp11_SPILL_256 <= Tspr11_2_V_0;
                       end 
                      
                  13'sd3300/*3300:xpc10*/:  begin 
                       xpc10 <= 13'sd3301/*3301:xpc10*/;
                       Tsf0SPILL12_256 <= 32'sd0;
                       end 
                      
                  13'sd3304/*3304:xpc10*/:  begin 
                       xpc10 <= 13'sd3305/*3305:xpc10*/;
                       Tsf0SPILL10_256 <= 32'sd0;
                       end 
                      
                  13'sd3317/*3317:xpc10*/:  begin 
                       xpc10 <= 13'sd3318/*3318:xpc10*/;
                       Tsf1SPILL10_256 <= 64'h_7fff_ffff_ffff_ffff;
                       end 
                      
                  13'sd3325/*3325:xpc10*/:  begin 
                       xpc10 <= 13'sd3326/*3326:xpc10*/;
                       Tsp15_SPILL_256 <= 64'sh1;
                       end 
                      
                  13'sd3329/*3329:xpc10*/:  begin 
                       xpc10 <= 13'sd3330/*3330:xpc10*/;
                       Tsf1SPILL10_256 <= $signed(64'sh_7ff0_0000_0000_0000+(Tsp15_SPILL_256<<32'sd63));
                       end 
                      
                  13'sd3333/*3333:xpc10*/:  begin 
                       xpc10 <= 13'sd3334/*3334:xpc10*/;
                       Tsp15_SPILL_256 <= 64'sh0;
                       end 
                      
                  13'sd3349/*3349:xpc10*/:  begin 
                       xpc10 <= 13'sd3350/*3350:xpc10*/;
                       Tsp18_SPILL_256 <= 64'sh1;
                       end 
                      
                  13'sd3353/*3353:xpc10*/:  begin 
                       xpc10 <= 13'sd3354/*3354:xpc10*/;
                       Tsf1SPILL10_256 <= $signed(64'sh0+(Tsp18_SPILL_256<<32'sd63));
                       end 
                      
                  13'sd3357/*3357:xpc10*/:  begin 
                       xpc10 <= 13'sd3358/*3358:xpc10*/;
                       Tsp18_SPILL_256 <= 64'sh0;
                       end 
                      
                  13'sd3361/*3361:xpc10*/:  begin 
                       xpc10 <= 13'sd3362/*3362:xpc10*/;
                       Tsco0_2_V_0 <= Tsfl1_24_V_6;
                       end 
                      
                  13'sd3362/*3362:xpc10*/:  begin 
                       xpc10 <= 13'sd3363/*3363:xpc10*/;
                       Tsco0_2_V_1 <= 8'h0;
                       end 
                      
                  13'sd3367/*3367:xpc10*/:  begin 
                       xpc10 <= 13'sd3368/*3368:xpc10*/;
                       Tsco0_2_V_1 <= 8'h20;
                       end 
                      
                  13'sd3371/*3371:xpc10*/:  begin 
                       xpc10 <= 13'sd3372/*3372:xpc10*/;
                       Tsco3_7_V_0 <= rtl_unsigned_bitextract6(64'h_ffff_ffff&Tsco0_2_V_0);
                       end 
                      
                  13'sd3372/*3372:xpc10*/:  begin 
                       xpc10 <= 13'sd3373/*3373:xpc10*/;
                       Tsco3_7_V_1 <= 8'h0;
                       end 
                      
                  13'sd3377/*3377:xpc10*/:  begin 
                       xpc10 <= 13'sd3378/*3378:xpc10*/;
                       Tsco3_7_V_1 <= 8'h10;
                       end 
                      
                  13'sd3378/*3378:xpc10*/:  begin 
                       xpc10 <= 13'sd3379/*3379:xpc10*/;
                       Tsco3_7_V_0 <= (Tsco3_7_V_0<<32'sd16);
                       end 
                      
                  13'sd3386/*3386:xpc10*/:  begin 
                       xpc10 <= 13'sd3387/*3387:xpc10*/;
                       Tsco3_7_V_1 <= rtl_unsigned_bitextract7(8'd8+Tsco3_7_V_1);
                       end 
                      
                  13'sd3387/*3387:xpc10*/:  begin 
                       xpc10 <= 13'sd3388/*3388:xpc10*/;
                       Tsco3_7_V_0 <= (Tsco3_7_V_0<<32'sd8);
                       end 
                      
                  13'sd3391/*3391:xpc10*/:  begin 
                       xpc10 <= 13'sd3392/*3392:xpc10*/;
                       Tsco3_7_V_1 <= rtl_unsigned_bitextract7(Tsco3_7_V_1+A_8_US_CC_SCALbx16_ARA0[$unsigned((Tsco3_7_V_0>>32'sd24))]
                      );

                       end 
                      
                  13'sd3392/*3392:xpc10*/:  begin 
                       xpc10 <= 13'sd3393/*3393:xpc10*/;
                       Tsco0_2_V_1 <= rtl_unsigned_bitextract7(Tsco0_2_V_1+Tsco3_7_V_1);
                       end 
                      
                  13'sd3393/*3393:xpc10*/:  begin 
                       xpc10 <= 13'sd3394/*3394:xpc10*/;
                       Tsno19_4_V_0 <= $unsigned(-32'sd11+rtl_sign_extend8(Tsco0_2_V_1));
                       end 
                      
                  13'sd3394/*3394:xpc10*/:  begin 
                       xpc10 <= 13'sd3395/*3395:xpc10*/;
                       Tsfl1_24_V_6 <= (Tsfl1_24_V_6<<(32'sd63&Tsno19_4_V_0));
                       end 
                      
                  13'sd3395/*3395:xpc10*/:  begin 
                       xpc10 <= 13'sd3396/*3396:xpc10*/;
                       Tsfl1_24_V_3 <= rtl_signed_bitextract0(rtl_sign_extend9(16'sd1)+(0-Tsno19_4_V_0));
                       end 
                      
                  13'sd3411/*3411:xpc10*/:  begin 
                       xpc10 <= 13'sd3412/*3412:xpc10*/;
                       Tsp22_SPILL_256 <= 64'sh1;
                       end 
                      
                  13'sd3415/*3415:xpc10*/:  begin 
                       xpc10 <= 13'sd3416/*3416:xpc10*/;
                       Tsf1SPILL10_256 <= $signed(64'sh0+(Tsp22_SPILL_256<<32'sd63));
                       end 
                      
                  13'sd3419/*3419:xpc10*/:  begin 
                       xpc10 <= 13'sd3420/*3420:xpc10*/;
                       Tsp22_SPILL_256 <= 64'sh0;
                       end 
                      
                  13'sd3423/*3423:xpc10*/:  begin 
                       xpc10 <= 13'sd3424/*3424:xpc10*/;
                       Tsco0_2_V_0 <= Tsfl1_24_V_7;
                       end 
                      
                  13'sd3424/*3424:xpc10*/:  begin 
                       xpc10 <= 13'sd3425/*3425:xpc10*/;
                       Tsco0_2_V_1 <= 8'h0;
                       end 
                      
                  13'sd3429/*3429:xpc10*/:  begin 
                       xpc10 <= 13'sd3430/*3430:xpc10*/;
                       Tsco0_2_V_1 <= 8'h20;
                       end 
                      
                  13'sd3433/*3433:xpc10*/:  begin 
                       xpc10 <= 13'sd3434/*3434:xpc10*/;
                       Tsco3_7_V_0 <= rtl_unsigned_bitextract6(64'h_ffff_ffff&Tsco0_2_V_0);
                       end 
                      
                  13'sd3434/*3434:xpc10*/:  begin 
                       xpc10 <= 13'sd3435/*3435:xpc10*/;
                       Tsco3_7_V_1 <= 8'h0;
                       end 
                      
                  13'sd3439/*3439:xpc10*/:  begin 
                       xpc10 <= 13'sd3440/*3440:xpc10*/;
                       Tsco3_7_V_1 <= 8'h10;
                       end 
                      
                  13'sd3440/*3440:xpc10*/:  begin 
                       xpc10 <= 13'sd3441/*3441:xpc10*/;
                       Tsco3_7_V_0 <= (Tsco3_7_V_0<<32'sd16);
                       end 
                      
                  13'sd3448/*3448:xpc10*/:  begin 
                       xpc10 <= 13'sd3449/*3449:xpc10*/;
                       Tsco3_7_V_1 <= rtl_unsigned_bitextract7(8'd8+Tsco3_7_V_1);
                       end 
                      
                  13'sd3449/*3449:xpc10*/:  begin 
                       xpc10 <= 13'sd3450/*3450:xpc10*/;
                       Tsco3_7_V_0 <= (Tsco3_7_V_0<<32'sd8);
                       end 
                      
                  13'sd3453/*3453:xpc10*/:  begin 
                       xpc10 <= 13'sd3454/*3454:xpc10*/;
                       Tsco3_7_V_1 <= rtl_unsigned_bitextract7(Tsco3_7_V_1+A_8_US_CC_SCALbx16_ARA0[$unsigned((Tsco3_7_V_0>>32'sd24))]
                      );

                       end 
                      
                  13'sd3454/*3454:xpc10*/:  begin 
                       xpc10 <= 13'sd3455/*3455:xpc10*/;
                       Tsco0_2_V_1 <= rtl_unsigned_bitextract7(Tsco0_2_V_1+Tsco3_7_V_1);
                       end 
                      
                  13'sd3455/*3455:xpc10*/:  begin 
                       xpc10 <= 13'sd3456/*3456:xpc10*/;
                       Tsno23_4_V_0 <= $unsigned(-32'sd11+rtl_sign_extend8(Tsco0_2_V_1));
                       end 
                      
                  13'sd3456/*3456:xpc10*/:  begin 
                       xpc10 <= 13'sd3457/*3457:xpc10*/;
                       Tsfl1_24_V_7 <= (Tsfl1_24_V_7<<(32'sd63&Tsno23_4_V_0));
                       end 
                      
                  13'sd3457/*3457:xpc10*/:  begin 
                       xpc10 <= 13'sd3458/*3458:xpc10*/;
                       Tsfl1_24_V_4 <= rtl_signed_bitextract0(rtl_sign_extend9(16'sd1)+(0-Tsno23_4_V_0));
                       end 
                      
                  13'sd3461/*3461:xpc10*/:  begin 
                       xpc10 <= 13'sd3462/*3462:xpc10*/;
                       Tsfl1_24_V_5 <= rtl_signed_bitextract0(-16'sd1023+Tsfl1_24_V_3+Tsfl1_24_V_4);
                       end 
                      
                  13'sd3462/*3462:xpc10*/:  begin 
                       xpc10 <= 13'sd3463/*3463:xpc10*/;
                       Tsfl1_24_V_6 <= ((64'sh10_0000_0000_0000|Tsfl1_24_V_6)<<32'sd10);
                       end 
                      
                  13'sd3463/*3463:xpc10*/:  begin 
                       xpc10 <= 13'sd3464/*3464:xpc10*/;
                       Tsfl1_24_V_7 <= ((64'sh10_0000_0000_0000|Tsfl1_24_V_7)<<32'sd11);
                       end 
                      
                  13'sd3464/*3464:xpc10*/:  begin 
                       xpc10 <= 13'sd3465/*3465:xpc10*/;
                       Tsmu24_24_V_1 <= rtl_unsigned_bitextract6(64'h_ffff_ffff&Tsfl1_24_V_6);
                       end 
                      
                  13'sd3465/*3465:xpc10*/:  begin 
                       xpc10 <= 13'sd3466/*3466:xpc10*/;
                       Tsmu24_24_V_0 <= rtl_unsigned_bitextract6((Tsfl1_24_V_6>>32'sd32));
                       end 
                      
                  13'sd3466/*3466:xpc10*/:  begin 
                       xpc10 <= 13'sd3467/*3467:xpc10*/;
                       Tsmu24_24_V_3 <= rtl_unsigned_bitextract6(64'h_ffff_ffff&Tsfl1_24_V_7);
                       end 
                      
                  13'sd3467/*3467:xpc10*/:  begin 
                       xpc10 <= 13'sd3468/*3468:xpc10*/;
                       Tsmu24_24_V_2 <= rtl_unsigned_bitextract6((Tsfl1_24_V_7>>32'sd32));
                       end 
                      
                  13'sd3468/*3468:xpc10*/:  begin 
                       xpc10 <= 13'sd3469/*3469:xpc10*/;
                       Tsmu24_24_V_7 <= rtl_unsigned_extend10(Tsmu24_24_V_1)*rtl_unsigned_extend10(Tsmu24_24_V_3);
                       end 
                      
                  13'sd3469/*3469:xpc10*/:  begin 
                       xpc10 <= 13'sd3470/*3470:xpc10*/;
                       Tsmu24_24_V_5 <= rtl_unsigned_extend10(Tsmu24_24_V_1)*rtl_unsigned_extend10(Tsmu24_24_V_2);
                       end 
                      
                  13'sd3470/*3470:xpc10*/:  begin 
                       xpc10 <= 13'sd3471/*3471:xpc10*/;
                       Tsmu24_24_V_6 <= rtl_unsigned_extend10(Tsmu24_24_V_0)*rtl_unsigned_extend10(Tsmu24_24_V_3);
                       end 
                      
                  13'sd3471/*3471:xpc10*/:  begin 
                       xpc10 <= 13'sd3472/*3472:xpc10*/;
                       Tsmu24_24_V_4 <= rtl_unsigned_extend10(Tsmu24_24_V_0)*rtl_unsigned_extend10(Tsmu24_24_V_2);
                       end 
                      
                  13'sd3472/*3472:xpc10*/:  begin 
                       xpc10 <= 13'sd3473/*3473:xpc10*/;
                       Tsmu24_24_V_5 <= Tsmu24_24_V_5+Tsmu24_24_V_6;
                       end 
                      
                  13'sd3482/*3482:xpc10*/:  begin 
                       xpc10 <= 13'sd3483/*3483:xpc10*/;
                       fastspilldup38 <= Tsmu24_24_V_4;
                       end 
                      
                  13'sd3483/*3483:xpc10*/:  begin 
                       xpc10 <= 13'sd3484/*3484:xpc10*/;
                       Tsm24_SPILL_264 <= fastspilldup38;
                       end 
                      
                  13'sd3484/*3484:xpc10*/:  begin 
                       xpc10 <= 13'sd3485/*3485:xpc10*/;
                       Tsm24_SPILL_257 <= fastspilldup38;
                       end 
                      
                  13'sd3489/*3489:xpc10*/:  begin 
                       xpc10 <= 13'sd3490/*3490:xpc10*/;
                       Tsm24_SPILL_259 <= 64'sh1;
                       end 
                      
                  13'sd3490/*3490:xpc10*/:  begin 
                       xpc10 <= 13'sd3491/*3491:xpc10*/;
                       Tsm24_SPILL_258 <= Tsm24_SPILL_257;
                       end 
                      
                  13'sd3494/*3494:xpc10*/:  begin 
                       xpc10 <= 13'sd3495/*3495:xpc10*/;
                       Tsmu24_24_V_4 <= Tsm24_SPILL_258+(Tsm24_SPILL_259<<32'sd32)+(Tsmu24_24_V_5>>32'sd32);
                       end 
                      
                  13'sd3495/*3495:xpc10*/:  begin 
                       xpc10 <= 13'sd3496/*3496:xpc10*/;
                       Tsmu24_24_V_5 <= (Tsmu24_24_V_5<<32'sd32);
                       end 
                      
                  13'sd3496/*3496:xpc10*/:  begin 
                       xpc10 <= 13'sd3497/*3497:xpc10*/;
                       Tsmu24_24_V_7 <= Tsmu24_24_V_7+Tsmu24_24_V_5;
                       end 
                      
                  13'sd3497/*3497:xpc10*/:  begin 
                       xpc10 <= 13'sd3498/*3498:xpc10*/;
                       fastspilldup40 <= Tsmu24_24_V_4;
                       end 
                      
                  13'sd3498/*3498:xpc10*/:  begin 
                       xpc10 <= 13'sd3499/*3499:xpc10*/;
                       Tsm24_SPILL_263 <= fastspilldup40;
                       end 
                      
                  13'sd3499/*3499:xpc10*/:  begin 
                       xpc10 <= 13'sd3500/*3500:xpc10*/;
                       Tsm24_SPILL_260 <= fastspilldup40;
                       end 
                      
                  13'sd3504/*3504:xpc10*/:  begin 
                       xpc10 <= 13'sd3505/*3505:xpc10*/;
                       Tsm24_SPILL_262 <= 64'sh1;
                       end 
                      
                  13'sd3505/*3505:xpc10*/:  begin 
                       xpc10 <= 13'sd3506/*3506:xpc10*/;
                       Tsm24_SPILL_261 <= Tsm24_SPILL_260;
                       end 
                      
                  13'sd3509/*3509:xpc10*/:  begin 
                       xpc10 <= 13'sd3510/*3510:xpc10*/;
                       Tsmu24_24_V_4 <= Tsm24_SPILL_262+Tsm24_SPILL_261;
                       end 
                      
                  13'sd3510/*3510:xpc10*/:  begin 
                       xpc10 <= 13'sd3511/*3511:xpc10*/;
                       Tsfl1_24_V_9 <= Tsmu24_24_V_7;
                       end 
                      
                  13'sd3511/*3511:xpc10*/:  begin 
                       xpc10 <= 13'sd3512/*3512:xpc10*/;
                       Tsfl1_24_V_8 <= Tsmu24_24_V_4;
                       end 
                      
                  13'sd3512/*3512:xpc10*/:  begin 
                       xpc10 <= 13'sd3513/*3513:xpc10*/;
                       fastspilldup42 <= Tsfl1_24_V_8;
                       end 
                      
                  13'sd3513/*3513:xpc10*/:  begin 
                       xpc10 <= 13'sd3514/*3514:xpc10*/;
                       Tsf1SPILL10_260 <= fastspilldup42;
                       end 
                      
                  13'sd3514/*3514:xpc10*/:  begin 
                       xpc10 <= 13'sd3515/*3515:xpc10*/;
                       Tsf1SPILL10_257 <= fastspilldup42;
                       end 
                      endcase
              if ((32'sd0/*0:USA74*/==(Tsro33_4_V_1<<(32'sd63&rtl_signed_bitextract0(Tsro33_4_V_0)))))  begin if ((13'sd2871/*2871:xpc10*/==
                  xpc10))  xpc10 <= 13'sd2882/*2882:xpc10*/;
                       end 
                   else if ((13'sd2871/*2871:xpc10*/==xpc10))  xpc10 <= 13'sd2872/*2872:xpc10*/;
                      
              case (xpc10)
                  13'sd2754/*2754:xpc10*/: if ((Tsro33_4_V_1+rtl_sign_extend1(Tsro33_4_V_5)<64'sh0))  xpc10 <= 13'sd2755/*2755:xpc10*/;
                       else  xpc10 <= 13'sd2794/*2794:xpc10*/;

                  13'sd2763/*2763:xpc10*/:  begin 
                       xpc10 <= 13'sd2764/*2764:xpc10*/;
                       Tsp13_SPILL_256 <= 64'sh1;
                       end 
                      
                  13'sd2767/*2767:xpc10*/:  begin 
                       xpc10 <= 13'sd2768/*2768:xpc10*/;
                       fastspilldup68 <= $signed(64'sh_7ff0_0000_0000_0000+(Tsp13_SPILL_256<<32'sd63));
                       end 
                      
                  13'sd2768/*2768:xpc10*/:  begin 
                       xpc10 <= 13'sd2769/*2769:xpc10*/;
                       Tsr33_SPILL_260 <= fastspilldup68;
                       end 
                      
                  13'sd2769/*2769:xpc10*/:  begin 
                       xpc10 <= 13'sd2770/*2770:xpc10*/;
                       Tsr33_SPILL_256 <= fastspilldup68;
                       end 
                      
                  13'sd2770/*2770:xpc10*/: if (!(!Tsro33_4_V_5))  xpc10 <= 13'sd2785/*2785:xpc10*/;
                       else  xpc10 <= 13'sd2771/*2771:xpc10*/;

                  13'sd2774/*2774:xpc10*/:  begin 
                       xpc10 <= 13'sd2775/*2775:xpc10*/;
                       Tsr33_SPILL_258 <= 64'sh1;
                       end 
                      
                  13'sd2775/*2775:xpc10*/:  begin 
                       xpc10 <= 13'sd2776/*2776:xpc10*/;
                       Tsr33_SPILL_257 <= Tsr33_SPILL_256;
                       end 
                      
                  13'sd2779/*2779:xpc10*/:  begin 
                       xpc10 <= 13'sd2780/*2780:xpc10*/;
                       Tsr33_SPILL_259 <= Tsr33_SPILL_257+(0-Tsr33_SPILL_258);
                       end 
                      
                  13'sd2783/*2783:xpc10*/:  begin 
                       xpc10 <= 13'sd2784/*2784:xpc10*/;
                       Tsf1SPILL12_256 <= Tsr33_SPILL_259;
                       end 
                      
                  13'sd2787/*2787:xpc10*/:  begin 
                       xpc10 <= 13'sd2788/*2788:xpc10*/;
                       Tsr33_SPILL_258 <= 64'sh0;
                       end 
                      
                  13'sd2788/*2788:xpc10*/:  begin 
                       xpc10 <= 13'sd2789/*2789:xpc10*/;
                       Tsr33_SPILL_257 <= Tsr33_SPILL_260;
                       end 
                      
                  13'sd2792/*2792:xpc10*/:  begin 
                       xpc10 <= 13'sd2793/*2793:xpc10*/;
                       Tsp13_SPILL_256 <= 64'sh0;
                       end 
                      
                  13'sd2796/*2796:xpc10*/: if ((Tsro33_4_V_0<32'sd0))  xpc10 <= 13'sd2797/*2797:xpc10*/;
                       else  xpc10 <= 13'sd2821/*2821:xpc10*/;

                  13'sd2801/*2801:xpc10*/: if (!(!rtl_signed_bitextract0((0-Tsro33_4_V_0))))  xpc10 <= 13'sd2862/*2862:xpc10*/;
                       else  xpc10 <= 13'sd2802/*2802:xpc10*/;

                  13'sd2805/*2805:xpc10*/:  begin 
                       xpc10 <= 13'sd2806/*2806:xpc10*/;
                       Tssh18_7_V_0 <= Tsro33_4_V_1;
                       end 
                      
                  13'sd2809/*2809:xpc10*/:  begin 
                       xpc10 <= 13'sd2810/*2810:xpc10*/;
                       Tsro33_4_V_1 <= Tssh18_7_V_0;
                       end 
                      
                  13'sd2810/*2810:xpc10*/:  begin 
                       xpc10 <= 13'sd2811/*2811:xpc10*/;
                       Tsro33_4_V_0 <= 16'sh0;
                       end 
                      
                  13'sd2811/*2811:xpc10*/:  begin 
                       xpc10 <= 13'sd2812/*2812:xpc10*/;
                       Tsro33_4_V_6 <= rtl_signed_bitextract2(64'sh3ff&Tsro33_4_V_1);
                       end 
                      
                  13'sd2831/*2831:xpc10*/:  begin 
                       xpc10 <= 13'sd2832/*2832:xpc10*/;
                       Tsro33_4_V_1 <= (Tsro33_4_V_1+rtl_sign_extend1(Tsro33_4_V_5)>>32'sd10);
                       end 
                      
                  13'sd2832/*2832:xpc10*/: if (32'sd1&(32'sd0/*0:USA76*/==(32'sd512^Tsro33_4_V_6)))  xpc10 <= 13'sd2833/*2833:xpc10*/;
                       else  xpc10 <= 13'sd2838/*2838:xpc10*/;

                  13'sd2836/*2836:xpc10*/:  begin 
                       xpc10 <= 13'sd2837/*2837:xpc10*/;
                       Tsro33_4_V_1 <= -64'sh2&Tsro33_4_V_1;
                       end 
                      
                  13'sd2844/*2844:xpc10*/:  begin 
                       xpc10 <= 13'sd2845/*2845:xpc10*/;
                       Tsro33_4_V_0 <= 16'sh0;
                       end 
                      
                  13'sd2852/*2852:xpc10*/:  begin 
                       xpc10 <= 13'sd2853/*2853:xpc10*/;
                       Tsp27_SPILL_256 <= 64'sh1;
                       end 
                      
                  13'sd2856/*2856:xpc10*/:  begin 
                       xpc10 <= 13'sd2857/*2857:xpc10*/;
                       Tsr33_SPILL_259 <= Tsro33_4_V_1+(Tsp27_SPILL_256<<32'sd63)+(rtl_sign_extend1(Tsro33_4_V_0)<<32'sd52);
                       end 
                      
                  13'sd2860/*2860:xpc10*/:  begin 
                       xpc10 <= 13'sd2861/*2861:xpc10*/;
                       Tsp27_SPILL_256 <= 64'sh0;
                       end 
                      
                  13'sd2864/*2864:xpc10*/: if ((rtl_signed_bitextract0((0-Tsro33_4_V_0))<32'sd64))  xpc10 <= 13'sd2865/*2865:xpc10*/;
                       else  xpc10 <= 13'sd2887/*2887:xpc10*/;

                  13'sd2868/*2868:xpc10*/:  begin 
                       xpc10 <= 13'sd2869/*2869:xpc10*/;
                       fastspilldup70 <= (Tsro33_4_V_1>>(32'sd63&rtl_signed_bitextract0((0-Tsro33_4_V_0))));
                       end 
                      
                  13'sd2869/*2869:xpc10*/:  begin 
                       xpc10 <= 13'sd2870/*2870:xpc10*/;
                       Tss18_SPILL_259 <= fastspilldup70;
                       end 
                      
                  13'sd2870/*2870:xpc10*/:  begin 
                       xpc10 <= 13'sd2871/*2871:xpc10*/;
                       Tss18_SPILL_256 <= fastspilldup70;
                       end 
                      endcase
              if ((Tsro33_4_V_0==32'sd2045/*2045:Tsro33.4_V_0*/))  begin if ((13'sd2750/*2750:xpc10*/==xpc10))  xpc10 <= 13'sd2751/*2751:xpc10*/;
                       end 
                   else if ((13'sd2750/*2750:xpc10*/==xpc10))  xpc10 <= 13'sd2794/*2794:xpc10*/;
                      
              case (xpc10)
                  13'sd2724/*2724:xpc10*/:  begin 
                       xpc10 <= 13'sd2725/*2725:xpc10*/;
                       Tsf1SPILL12_259 <= 64'sh1;
                       end 
                      
                  13'sd2725/*2725:xpc10*/:  begin 
                       xpc10 <= 13'sd2726/*2726:xpc10*/;
                       Tsf1SPILL12_258 <= Tsf1SPILL12_257;
                       end 
                      
                  13'sd2729/*2729:xpc10*/:  begin 
                       xpc10 <= 13'sd2730/*2730:xpc10*/;
                       Tsfl1_35_V_8 <= Tsf1SPILL12_259|Tsf1SPILL12_258;
                       end 
                      
                  13'sd2733/*2733:xpc10*/:  begin 
                       xpc10 <= 13'sd2734/*2734:xpc10*/;
                       Tsro33_4_V_0 <= rtl_signed_bitextract0(Tsfl1_35_V_5);
                       end 
                      
                  13'sd2734/*2734:xpc10*/:  begin 
                       xpc10 <= 13'sd2735/*2735:xpc10*/;
                       Tsro33_4_V_1 <= Tsfl1_35_V_8;
                       end 
                      
                  13'sd2737/*2737:xpc10*/:  begin 
                       xpc10 <= 13'sd2738/*2738:xpc10*/;
                       Tsro33_4_V_5 <= 16'sh200;
                       end 
                      
                  13'sd2741/*2741:xpc10*/:  begin 
                       xpc10 <= 13'sd2742/*2742:xpc10*/;
                       Tsro33_4_V_6 <= rtl_signed_bitextract2(64'sh3ff&Tsro33_4_V_1);
                       end 
                      
                  13'sd2742/*2742:xpc10*/: if ((Tsro33_4_V_0<32'sd2045))  xpc10 <= 13'sd2821/*2821:xpc10*/;
                       else  xpc10 <= 13'sd2743/*2743:xpc10*/;

                  13'sd2746/*2746:xpc10*/: if ((32'sd2045<Tsro33_4_V_0))  xpc10 <= 13'sd2756/*2756:xpc10*/;
                       else  xpc10 <= 13'sd2747/*2747:xpc10*/;
              endcase
              if ((Tsfl1_35_V_10==32'sd0/*0:Tsfl1.35_V_10*/))  begin if ((13'sd2720/*2720:xpc10*/==xpc10))  xpc10 <= 13'sd2903/*2903:xpc10*/;
                       end 
                   else if ((13'sd2720/*2720:xpc10*/==xpc10))  xpc10 <= 13'sd2721/*2721:xpc10*/;
                      
              case (xpc10)
                  13'sd2414/*2414:xpc10*/:  begin 
                       xpc10 <= 13'sd2415/*2415:xpc10*/;
                       Tsf0SPILL12_256 <= rtl_sign_extend3((32'sd0/*0:USA72*/==(32'sd0/*0:USA70*/==(64'sh7_ffff_ffff_ffff&Tspr10_2_V_1
                      ))));

                       end 
                      
                  13'sd2418/*2418:xpc10*/:  begin 
                       xpc10 <= 13'sd2419/*2419:xpc10*/;
                       Tspr10_2_V_4 <= rtl_unsigned_bitextract4(Tsf0SPILL12_256);
                       end 
                      
                  13'sd2419/*2419:xpc10*/:  begin 
                       xpc10 <= 13'sd2420/*2420:xpc10*/;
                       Tspr10_2_V_0 <= 64'sh8_0000_0000_0000|Tspr10_2_V_0;
                       end 
                      
                  13'sd2420/*2420:xpc10*/:  begin 
                       xpc10 <= 13'sd2421/*2421:xpc10*/;
                       Tspr10_2_V_1 <= 64'sh8_0000_0000_0000|Tspr10_2_V_1;
                       end 
                      
                  13'sd2421/*2421:xpc10*/:  begin 
                      if (Tspr10_2_V_2 || Tspr10_2_V_4)  begin if (Tspr10_2_V_2 || Tspr10_2_V_4)  xpc10 <= 13'sd2422/*2422:xpc10*/;
                               end 
                          if (!Tspr10_2_V_2 && !Tspr10_2_V_4)  xpc10 <= 13'sd2427/*2427:xpc10*/;
                           end 
                      
                  13'sd2429/*2429:xpc10*/: if (Tspr10_2_V_4)  xpc10 <= 13'sd2430/*2430:xpc10*/;
                       else  xpc10 <= 13'sd2439/*2439:xpc10*/;

                  13'sd2433/*2433:xpc10*/:  begin 
                       xpc10 <= 13'sd2434/*2434:xpc10*/;
                       Tsp10_SPILL_256 <= Tspr10_2_V_1;
                       end 
                      
                  13'sd2437/*2437:xpc10*/:  begin 
                       xpc10 <= 13'sd2438/*2438:xpc10*/;
                       Tsf1SPILL12_256 <= Tsp10_SPILL_256;
                       end 
                      
                  13'sd2441/*2441:xpc10*/: if (Tspr10_2_V_2)  xpc10 <= 13'sd2442/*2442:xpc10*/;
                       else  xpc10 <= 13'sd2447/*2447:xpc10*/;

                  13'sd2445/*2445:xpc10*/:  begin 
                       xpc10 <= 13'sd2446/*2446:xpc10*/;
                       Tsp10_SPILL_256 <= Tspr10_2_V_0;
                       end 
                      
                  13'sd2449/*2449:xpc10*/: if (Tspr10_2_V_3)  xpc10 <= 13'sd2450/*2450:xpc10*/;
                       else  xpc10 <= 13'sd2455/*2455:xpc10*/;

                  13'sd2453/*2453:xpc10*/:  begin 
                       xpc10 <= 13'sd2454/*2454:xpc10*/;
                       Tsp10_SPILL_256 <= Tspr10_2_V_1;
                       end 
                      
                  13'sd2457/*2457:xpc10*/:  begin 
                       xpc10 <= 13'sd2458/*2458:xpc10*/;
                       Tsp10_SPILL_256 <= Tspr10_2_V_0;
                       end 
                      
                  13'sd2461/*2461:xpc10*/:  begin 
                       xpc10 <= 13'sd2462/*2462:xpc10*/;
                       Tsf0SPILL12_256 <= 32'sd0;
                       end 
                      
                  13'sd2465/*2465:xpc10*/:  begin 
                       xpc10 <= 13'sd2466/*2466:xpc10*/;
                       Tsf0SPILL10_256 <= 32'sd0;
                       end 
                      
                  13'sd2473/*2473:xpc10*/:  begin 
                       xpc10 <= 13'sd2474/*2474:xpc10*/;
                       Tsp11SPILL10_256 <= 64'sh1;
                       end 
                      
                  13'sd2477/*2477:xpc10*/:  begin 
                       xpc10 <= 13'sd2478/*2478:xpc10*/;
                       Tsf1SPILL12_256 <= $signed(64'sh0+(Tsp11SPILL10_256<<32'sd63));
                       end 
                      
                  13'sd2481/*2481:xpc10*/:  begin 
                       xpc10 <= 13'sd2482/*2482:xpc10*/;
                       Tsp11SPILL10_256 <= 64'sh0;
                       end 
                      
                  13'sd2485/*2485:xpc10*/: if (!(!Tsfl1_35_V_4))  xpc10 <= 13'sd2559/*2559:xpc10*/;
                       else  xpc10 <= 13'sd2486/*2486:xpc10*/;

                  13'sd2502/*2502:xpc10*/:  begin 
                       xpc10 <= 13'sd2503/*2503:xpc10*/;
                       Tsf1SPILL12_256 <= 64'h_7fff_ffff_ffff_ffff;
                       end 
                      
                  13'sd2511/*2511:xpc10*/:  begin 
                       xpc10 <= 13'sd2512/*2512:xpc10*/;
                       Tsp17_SPILL_256 <= 64'sh1;
                       end 
                      
                  13'sd2515/*2515:xpc10*/:  begin 
                       xpc10 <= 13'sd2516/*2516:xpc10*/;
                       Tsf1SPILL12_256 <= $signed(64'sh_7ff0_0000_0000_0000+(Tsp17_SPILL_256<<32'sd63));
                       end 
                      
                  13'sd2519/*2519:xpc10*/:  begin 
                       xpc10 <= 13'sd2520/*2520:xpc10*/;
                       Tsp17_SPILL_256 <= 64'sh0;
                       end 
                      
                  13'sd2523/*2523:xpc10*/:  begin 
                       xpc10 <= 13'sd2524/*2524:xpc10*/;
                       Tsco0_2_V_0 <= Tsfl1_35_V_7;
                       end 
                      
                  13'sd2524/*2524:xpc10*/:  begin 
                       xpc10 <= 13'sd2525/*2525:xpc10*/;
                       Tsco0_2_V_1 <= 8'h0;
                       end 
                      
                  13'sd2529/*2529:xpc10*/:  begin 
                       xpc10 <= 13'sd2530/*2530:xpc10*/;
                       Tsco0_2_V_1 <= 8'h20;
                       end 
                      
                  13'sd2533/*2533:xpc10*/:  begin 
                       xpc10 <= 13'sd2534/*2534:xpc10*/;
                       Tsco3_7_V_0 <= rtl_unsigned_bitextract6(64'h_ffff_ffff&Tsco0_2_V_0);
                       end 
                      
                  13'sd2534/*2534:xpc10*/:  begin 
                       xpc10 <= 13'sd2535/*2535:xpc10*/;
                       Tsco3_7_V_1 <= 8'h0;
                       end 
                      
                  13'sd2539/*2539:xpc10*/:  begin 
                       xpc10 <= 13'sd2540/*2540:xpc10*/;
                       Tsco3_7_V_1 <= 8'h10;
                       end 
                      
                  13'sd2540/*2540:xpc10*/:  begin 
                       xpc10 <= 13'sd2541/*2541:xpc10*/;
                       Tsco3_7_V_0 <= (Tsco3_7_V_0<<32'sd16);
                       end 
                      
                  13'sd2548/*2548:xpc10*/:  begin 
                       xpc10 <= 13'sd2549/*2549:xpc10*/;
                       Tsco3_7_V_1 <= rtl_unsigned_bitextract7(8'd8+Tsco3_7_V_1);
                       end 
                      
                  13'sd2549/*2549:xpc10*/:  begin 
                       xpc10 <= 13'sd2550/*2550:xpc10*/;
                       Tsco3_7_V_0 <= (Tsco3_7_V_0<<32'sd8);
                       end 
                      
                  13'sd2553/*2553:xpc10*/:  begin 
                       xpc10 <= 13'sd2554/*2554:xpc10*/;
                       Tsco3_7_V_1 <= rtl_unsigned_bitextract7(Tsco3_7_V_1+A_8_US_CC_SCALbx16_ARA0[$unsigned((Tsco3_7_V_0>>32'sd24))]
                      );

                       end 
                      
                  13'sd2554/*2554:xpc10*/:  begin 
                       xpc10 <= 13'sd2555/*2555:xpc10*/;
                       Tsco0_2_V_1 <= rtl_unsigned_bitextract7(Tsco0_2_V_1+Tsco3_7_V_1);
                       end 
                      
                  13'sd2555/*2555:xpc10*/:  begin 
                       xpc10 <= 13'sd2556/*2556:xpc10*/;
                       Tsno18_4_V_0 <= $unsigned(-32'sd11+rtl_sign_extend8(Tsco0_2_V_1));
                       end 
                      
                  13'sd2556/*2556:xpc10*/:  begin 
                       xpc10 <= 13'sd2557/*2557:xpc10*/;
                       Tsfl1_35_V_7 <= (Tsfl1_35_V_7<<(32'sd63&Tsno18_4_V_0));
                       end 
                      
                  13'sd2557/*2557:xpc10*/:  begin 
                       xpc10 <= 13'sd2558/*2558:xpc10*/;
                       Tsfl1_35_V_4 <= rtl_signed_bitextract0(rtl_sign_extend9(16'sd1)+(0-Tsno18_4_V_0));
                       end 
                      
                  13'sd2573/*2573:xpc10*/:  begin 
                       xpc10 <= 13'sd2574/*2574:xpc10*/;
                       Tsp21_SPILL_256 <= 64'sh1;
                       end 
                      
                  13'sd2577/*2577:xpc10*/:  begin 
                       xpc10 <= 13'sd2578/*2578:xpc10*/;
                       Tsf1SPILL12_256 <= $signed(64'sh0+(Tsp21_SPILL_256<<32'sd63));
                       end 
                      
                  13'sd2581/*2581:xpc10*/:  begin 
                       xpc10 <= 13'sd2582/*2582:xpc10*/;
                       Tsp21_SPILL_256 <= 64'sh0;
                       end 
                      
                  13'sd2585/*2585:xpc10*/:  begin 
                       xpc10 <= 13'sd2586/*2586:xpc10*/;
                       Tsco0_2_V_0 <= Tsfl1_35_V_6;
                       end 
                      
                  13'sd2586/*2586:xpc10*/:  begin 
                       xpc10 <= 13'sd2587/*2587:xpc10*/;
                       Tsco0_2_V_1 <= 8'h0;
                       end 
                      
                  13'sd2591/*2591:xpc10*/:  begin 
                       xpc10 <= 13'sd2592/*2592:xpc10*/;
                       Tsco0_2_V_1 <= 8'h20;
                       end 
                      
                  13'sd2595/*2595:xpc10*/:  begin 
                       xpc10 <= 13'sd2596/*2596:xpc10*/;
                       Tsco3_7_V_0 <= rtl_unsigned_bitextract6(64'h_ffff_ffff&Tsco0_2_V_0);
                       end 
                      
                  13'sd2596/*2596:xpc10*/:  begin 
                       xpc10 <= 13'sd2597/*2597:xpc10*/;
                       Tsco3_7_V_1 <= 8'h0;
                       end 
                      
                  13'sd2601/*2601:xpc10*/:  begin 
                       xpc10 <= 13'sd2602/*2602:xpc10*/;
                       Tsco3_7_V_1 <= 8'h10;
                       end 
                      
                  13'sd2602/*2602:xpc10*/:  begin 
                       xpc10 <= 13'sd2603/*2603:xpc10*/;
                       Tsco3_7_V_0 <= (Tsco3_7_V_0<<32'sd16);
                       end 
                      
                  13'sd2610/*2610:xpc10*/:  begin 
                       xpc10 <= 13'sd2611/*2611:xpc10*/;
                       Tsco3_7_V_1 <= rtl_unsigned_bitextract7(8'd8+Tsco3_7_V_1);
                       end 
                      
                  13'sd2611/*2611:xpc10*/:  begin 
                       xpc10 <= 13'sd2612/*2612:xpc10*/;
                       Tsco3_7_V_0 <= (Tsco3_7_V_0<<32'sd8);
                       end 
                      
                  13'sd2615/*2615:xpc10*/:  begin 
                       xpc10 <= 13'sd2616/*2616:xpc10*/;
                       Tsco3_7_V_1 <= rtl_unsigned_bitextract7(Tsco3_7_V_1+A_8_US_CC_SCALbx16_ARA0[$unsigned((Tsco3_7_V_0>>32'sd24))]
                      );

                       end 
                      
                  13'sd2616/*2616:xpc10*/:  begin 
                       xpc10 <= 13'sd2617/*2617:xpc10*/;
                       Tsco0_2_V_1 <= rtl_unsigned_bitextract7(Tsco0_2_V_1+Tsco3_7_V_1);
                       end 
                      
                  13'sd2617/*2617:xpc10*/:  begin 
                       xpc10 <= 13'sd2618/*2618:xpc10*/;
                       Tsno22_4_V_0 <= $unsigned(-32'sd11+rtl_sign_extend8(Tsco0_2_V_1));
                       end 
                      
                  13'sd2618/*2618:xpc10*/:  begin 
                       xpc10 <= 13'sd2619/*2619:xpc10*/;
                       Tsfl1_35_V_6 <= (Tsfl1_35_V_6<<(32'sd63&Tsno22_4_V_0));
                       end 
                      
                  13'sd2619/*2619:xpc10*/:  begin 
                       xpc10 <= 13'sd2620/*2620:xpc10*/;
                       Tsfl1_35_V_3 <= rtl_signed_bitextract0(rtl_sign_extend9(16'sd1)+(0-Tsno22_4_V_0));
                       end 
                      
                  13'sd2623/*2623:xpc10*/:  begin 
                       xpc10 <= 13'sd2624/*2624:xpc10*/;
                       Tsfl1_35_V_5 <= rtl_signed_bitextract0(rtl_sign_extend9(16'sd1021)+rtl_sign_extend9(Tsfl1_35_V_3)+(0-Tsfl1_35_V_4
                      ));

                       end 
                      
                  13'sd2624/*2624:xpc10*/:  begin 
                       xpc10 <= 13'sd2625/*2625:xpc10*/;
                       Tsfl1_35_V_6 <= ((64'sh10_0000_0000_0000|Tsfl1_35_V_6)<<32'sd10);
                       end 
                      
                  13'sd2625/*2625:xpc10*/:  begin 
                       xpc10 <= 13'sd2626/*2626:xpc10*/;
                       Tsfl1_35_V_7 <= ((64'sh10_0000_0000_0000|Tsfl1_35_V_7)<<32'sd11);
                       end 
                      
                  13'sd2626/*2626:xpc10*/: if ((Tsfl1_35_V_6+Tsfl1_35_V_6<Tsfl1_35_V_7))  xpc10 <= 13'sd2633/*2633:xpc10*/;
                       else  xpc10 <= 13'sd2627/*2627:xpc10*/;

                  13'sd2630/*2630:xpc10*/:  begin 
                       xpc10 <= 13'sd2631/*2631:xpc10*/;
                       Tsfl1_35_V_6 <= (Tsfl1_35_V_6>>32'sd1);
                       end 
                      
                  13'sd2631/*2631:xpc10*/:  begin 
                       xpc10 <= 13'sd2632/*2632:xpc10*/;
                       Tsfl1_35_V_5 <= rtl_signed_bitextract0(16'sd1+Tsfl1_35_V_5);
                       end 
                      
                  13'sd2635/*2635:xpc10*/: if ((Tsfl1_35_V_6<Tsfl1_35_V_7))  xpc10 <= 13'sd2951/*2951:xpc10*/;
                       else  xpc10 <= 13'sd2636/*2636:xpc10*/;

                  13'sd2639/*2639:xpc10*/:  begin 
                       xpc10 <= 13'sd2640/*2640:xpc10*/;
                       Tse25_SPILL_256 <= 64'h_ffff_ffff_ffff_ffff;
                       end 
                      
                  13'sd2643/*2643:xpc10*/:  begin 
                       xpc10 <= 13'sd2644/*2644:xpc10*/;
                       Tsfl1_35_V_8 <= Tse25_SPILL_256;
                       end 
                      
                  13'sd2644/*2644:xpc10*/: if ((64'sh2<(64'sh1ff&Tsfl1_35_V_8)))  xpc10 <= 13'sd2731/*2731:xpc10*/;
                       else  xpc10 <= 13'sd2645/*2645:xpc10*/;

                  13'sd2648/*2648:xpc10*/:  begin 
                       xpc10 <= 13'sd2649/*2649:xpc10*/;
                       Tsmu26_4_V_1 <= rtl_unsigned_bitextract6(64'h_ffff_ffff&Tsfl1_35_V_7);
                       end 
                      
                  13'sd2649/*2649:xpc10*/:  begin 
                       xpc10 <= 13'sd2650/*2650:xpc10*/;
                       Tsmu26_4_V_0 <= rtl_unsigned_bitextract6((Tsfl1_35_V_7>>32'sd32));
                       end 
                      
                  13'sd2650/*2650:xpc10*/:  begin 
                       xpc10 <= 13'sd2651/*2651:xpc10*/;
                       Tsmu26_4_V_3 <= rtl_unsigned_bitextract6(64'h_ffff_ffff&Tsfl1_35_V_8);
                       end 
                      
                  13'sd2651/*2651:xpc10*/:  begin 
                       xpc10 <= 13'sd2652/*2652:xpc10*/;
                       Tsmu26_4_V_2 <= rtl_unsigned_bitextract6((Tsfl1_35_V_8>>32'sd32));
                       end 
                      
                  13'sd2652/*2652:xpc10*/:  begin 
                       xpc10 <= 13'sd2653/*2653:xpc10*/;
                       Tsmu26_4_V_7 <= rtl_unsigned_extend10(Tsmu26_4_V_1)*rtl_unsigned_extend10(Tsmu26_4_V_3);
                       end 
                      
                  13'sd2653/*2653:xpc10*/:  begin 
                       xpc10 <= 13'sd2654/*2654:xpc10*/;
                       Tsmu26_4_V_5 <= rtl_unsigned_extend10(Tsmu26_4_V_1)*rtl_unsigned_extend10(Tsmu26_4_V_2);
                       end 
                      
                  13'sd2654/*2654:xpc10*/:  begin 
                       xpc10 <= 13'sd2655/*2655:xpc10*/;
                       Tsmu26_4_V_6 <= rtl_unsigned_extend10(Tsmu26_4_V_0)*rtl_unsigned_extend10(Tsmu26_4_V_3);
                       end 
                      
                  13'sd2655/*2655:xpc10*/:  begin 
                       xpc10 <= 13'sd2656/*2656:xpc10*/;
                       Tsmu26_4_V_4 <= rtl_unsigned_extend10(Tsmu26_4_V_0)*rtl_unsigned_extend10(Tsmu26_4_V_2);
                       end 
                      
                  13'sd2656/*2656:xpc10*/:  begin 
                       xpc10 <= 13'sd2657/*2657:xpc10*/;
                       Tsmu26_4_V_5 <= Tsmu26_4_V_5+Tsmu26_4_V_6;
                       end 
                      
                  13'sd2666/*2666:xpc10*/:  begin 
                       xpc10 <= 13'sd2667/*2667:xpc10*/;
                       fastspilldup58 <= Tsmu26_4_V_4;
                       end 
                      
                  13'sd2667/*2667:xpc10*/:  begin 
                       xpc10 <= 13'sd2668/*2668:xpc10*/;
                       Tsm26_SPILL_264 <= fastspilldup58;
                       end 
                      
                  13'sd2668/*2668:xpc10*/:  begin 
                       xpc10 <= 13'sd2669/*2669:xpc10*/;
                       Tsm26_SPILL_257 <= fastspilldup58;
                       end 
                      
                  13'sd2673/*2673:xpc10*/:  begin 
                       xpc10 <= 13'sd2674/*2674:xpc10*/;
                       Tsm26_SPILL_259 <= 64'sh1;
                       end 
                      
                  13'sd2674/*2674:xpc10*/:  begin 
                       xpc10 <= 13'sd2675/*2675:xpc10*/;
                       Tsm26_SPILL_258 <= Tsm26_SPILL_257;
                       end 
                      
                  13'sd2678/*2678:xpc10*/:  begin 
                       xpc10 <= 13'sd2679/*2679:xpc10*/;
                       Tsmu26_4_V_4 <= Tsm26_SPILL_258+(Tsm26_SPILL_259<<32'sd32)+(Tsmu26_4_V_5>>32'sd32);
                       end 
                      
                  13'sd2679/*2679:xpc10*/:  begin 
                       xpc10 <= 13'sd2680/*2680:xpc10*/;
                       Tsmu26_4_V_5 <= (Tsmu26_4_V_5<<32'sd32);
                       end 
                      
                  13'sd2680/*2680:xpc10*/:  begin 
                       xpc10 <= 13'sd2681/*2681:xpc10*/;
                       Tsmu26_4_V_7 <= Tsmu26_4_V_7+Tsmu26_4_V_5;
                       end 
                      
                  13'sd2681/*2681:xpc10*/:  begin 
                       xpc10 <= 13'sd2682/*2682:xpc10*/;
                       fastspilldup60 <= Tsmu26_4_V_4;
                       end 
                      
                  13'sd2682/*2682:xpc10*/:  begin 
                       xpc10 <= 13'sd2683/*2683:xpc10*/;
                       Tsm26_SPILL_263 <= fastspilldup60;
                       end 
                      
                  13'sd2683/*2683:xpc10*/:  begin 
                       xpc10 <= 13'sd2684/*2684:xpc10*/;
                       Tsm26_SPILL_260 <= fastspilldup60;
                       end 
                      
                  13'sd2684/*2684:xpc10*/: if ((Tsmu26_4_V_7<Tsmu26_4_V_5))  xpc10 <= 13'sd2685/*2685:xpc10*/;
                       else  xpc10 <= 13'sd2937/*2937:xpc10*/;

                  13'sd2688/*2688:xpc10*/:  begin 
                       xpc10 <= 13'sd2689/*2689:xpc10*/;
                       Tsm26_SPILL_262 <= 64'sh1;
                       end 
                      
                  13'sd2689/*2689:xpc10*/:  begin 
                       xpc10 <= 13'sd2690/*2690:xpc10*/;
                       Tsm26_SPILL_261 <= Tsm26_SPILL_260;
                       end 
                      
                  13'sd2693/*2693:xpc10*/:  begin 
                       xpc10 <= 13'sd2694/*2694:xpc10*/;
                       Tsmu26_4_V_4 <= Tsm26_SPILL_262+Tsm26_SPILL_261;
                       end 
                      
                  13'sd2694/*2694:xpc10*/:  begin 
                       xpc10 <= 13'sd2695/*2695:xpc10*/;
                       Tsfl1_35_V_12 <= Tsmu26_4_V_7;
                       end 
                      
                  13'sd2695/*2695:xpc10*/:  begin 
                       xpc10 <= 13'sd2696/*2696:xpc10*/;
                       Tsfl1_35_V_11 <= Tsmu26_4_V_4;
                       end 
                      
                  13'sd2696/*2696:xpc10*/:  begin 
                       xpc10 <= 13'sd2697/*2697:xpc10*/;
                       Tsfl1_35_V_10 <= 64'sh0+(0-Tsfl1_35_V_12);
                       end 
                      
                  13'sd2697/*2697:xpc10*/:  begin 
                       xpc10 <= 13'sd2698/*2698:xpc10*/;
                       fastspilldup62 <= Tsfl1_35_V_6+(0-Tsfl1_35_V_11);
                       end 
                      
                  13'sd2698/*2698:xpc10*/:  begin 
                       xpc10 <= 13'sd2699/*2699:xpc10*/;
                       Tss26_SPILL_262 <= fastspilldup62;
                       end 
                      
                  13'sd2699/*2699:xpc10*/:  begin 
                       xpc10 <= 13'sd2700/*2700:xpc10*/;
                       Tss26_SPILL_257 <= fastspilldup62;
                       end 
                      
                  13'sd2700/*2700:xpc10*/: if ((64'sh0<Tsfl1_35_V_12))  xpc10 <= 13'sd2701/*2701:xpc10*/;
                       else  xpc10 <= 13'sd2932/*2932:xpc10*/;

                  13'sd2704/*2704:xpc10*/:  begin 
                       xpc10 <= 13'sd2705/*2705:xpc10*/;
                       Tss26_SPILL_260 <= 64'sh1;
                       end 
                      
                  13'sd2705/*2705:xpc10*/:  begin 
                       xpc10 <= 13'sd2706/*2706:xpc10*/;
                       Tss26_SPILL_259 <= Tss26_SPILL_257;
                       end 
                      
                  13'sd2709/*2709:xpc10*/:  begin 
                       xpc10 <= 13'sd2710/*2710:xpc10*/;
                       Tsfl1_35_V_9 <= Tss26_SPILL_259+(0-Tss26_SPILL_260);
                       end 
                      
                  13'sd2713/*2713:xpc10*/: if ((Tsfl1_35_V_9<64'sh0))  xpc10 <= 13'sd2908/*2908:xpc10*/;
                       else  xpc10 <= 13'sd2714/*2714:xpc10*/;

                  13'sd2717/*2717:xpc10*/:  begin 
                       xpc10 <= 13'sd2718/*2718:xpc10*/;
                       fastspilldup66 <= Tsfl1_35_V_8;
                       end 
                      
                  13'sd2718/*2718:xpc10*/:  begin 
                       xpc10 <= 13'sd2719/*2719:xpc10*/;
                       Tsf1SPILL12_260 <= fastspilldup66;
                       end 
                      
                  13'sd2719/*2719:xpc10*/:  begin 
                       xpc10 <= 13'sd2720/*2720:xpc10*/;
                       Tsf1SPILL12_257 <= fastspilldup66;
                       end 
                      endcase
              if ((32'sd4094/*4094:USA68*/==(64'shfff&(Tspr10_2_V_1>>32'sd51))))  begin if ((13'sd2410/*2410:xpc10*/==xpc10))  xpc10 <= 13'sd2411
                      /*2411:xpc10*/;

                       end 
                   else if ((13'sd2410/*2410:xpc10*/==xpc10))  xpc10 <= 13'sd2459/*2459:xpc10*/;
                      
              case (xpc10)
                  13'sd2404/*2404:xpc10*/:  begin 
                       xpc10 <= 13'sd2405/*2405:xpc10*/;
                       Tsf0SPILL10_256 <= rtl_sign_extend3((32'sd0/*0:USA66*/==(32'sd0/*0:USA64*/==(64'sh7_ffff_ffff_ffff&Tspr10_2_V_0
                      ))));

                       end 
                      
                  13'sd2408/*2408:xpc10*/:  begin 
                       xpc10 <= 13'sd2409/*2409:xpc10*/;
                       Tspr10_2_V_2 <= rtl_unsigned_bitextract4(Tsf0SPILL10_256);
                       end 
                      
                  13'sd2409/*2409:xpc10*/:  begin 
                       xpc10 <= 13'sd2410/*2410:xpc10*/;
                       Tspr10_2_V_3 <= (32'sd0<rtl_sign_extend5(54'sd9007199254740992)+(Tspr10_2_V_1<<32'sd1));
                       end 
                      endcase
              if ((32'sd4094/*4094:USA62*/==(64'shfff&(Tspr10_2_V_0>>32'sd51))))  begin if ((13'sd2400/*2400:xpc10*/==xpc10))  xpc10 <= 13'sd2401
                      /*2401:xpc10*/;

                       end 
                   else if ((13'sd2400/*2400:xpc10*/==xpc10))  xpc10 <= 13'sd2463/*2463:xpc10*/;
                      
              case (xpc10)
                  13'sd2314/*2314:xpc10*/:  begin 
                       xpc10 <= 13'sd2315/*2315:xpc10*/;
                       Tsf0SPILL12_256 <= rtl_sign_extend3((32'sd0/*0:USA60*/==(32'sd0/*0:USA58*/==(64'sh7_ffff_ffff_ffff&Tspr5_2_V_1
                      ))));

                       end 
                      
                  13'sd2318/*2318:xpc10*/:  begin 
                       xpc10 <= 13'sd2319/*2319:xpc10*/;
                       Tspr5_2_V_4 <= rtl_unsigned_bitextract4(Tsf0SPILL12_256);
                       end 
                      
                  13'sd2319/*2319:xpc10*/:  begin 
                       xpc10 <= 13'sd2320/*2320:xpc10*/;
                       Tspr5_2_V_0 <= 64'sh8_0000_0000_0000|Tspr5_2_V_0;
                       end 
                      
                  13'sd2320/*2320:xpc10*/:  begin 
                       xpc10 <= 13'sd2321/*2321:xpc10*/;
                       Tspr5_2_V_1 <= 64'sh8_0000_0000_0000|Tspr5_2_V_1;
                       end 
                      
                  13'sd2321/*2321:xpc10*/:  begin 
                      if (Tspr5_2_V_2 || Tspr5_2_V_4)  begin if (Tspr5_2_V_2 || Tspr5_2_V_4)  xpc10 <= 13'sd2322/*2322:xpc10*/;
                               end 
                          if (!Tspr5_2_V_2 && !Tspr5_2_V_4)  xpc10 <= 13'sd2327/*2327:xpc10*/;
                           end 
                      
                  13'sd2329/*2329:xpc10*/: if (Tspr5_2_V_4)  xpc10 <= 13'sd2330/*2330:xpc10*/;
                       else  xpc10 <= 13'sd2339/*2339:xpc10*/;

                  13'sd2333/*2333:xpc10*/:  begin 
                       xpc10 <= 13'sd2334/*2334:xpc10*/;
                       Tsp5SPILL10_256 <= Tspr5_2_V_1;
                       end 
                      
                  13'sd2337/*2337:xpc10*/:  begin 
                       xpc10 <= 13'sd2338/*2338:xpc10*/;
                       Tsf1SPILL12_256 <= Tsp5SPILL10_256;
                       end 
                      
                  13'sd2341/*2341:xpc10*/: if (Tspr5_2_V_2)  xpc10 <= 13'sd2342/*2342:xpc10*/;
                       else  xpc10 <= 13'sd2347/*2347:xpc10*/;

                  13'sd2345/*2345:xpc10*/:  begin 
                       xpc10 <= 13'sd2346/*2346:xpc10*/;
                       Tsp5SPILL10_256 <= Tspr5_2_V_0;
                       end 
                      
                  13'sd2349/*2349:xpc10*/: if (Tspr5_2_V_3)  xpc10 <= 13'sd2350/*2350:xpc10*/;
                       else  xpc10 <= 13'sd2355/*2355:xpc10*/;

                  13'sd2353/*2353:xpc10*/:  begin 
                       xpc10 <= 13'sd2354/*2354:xpc10*/;
                       Tsp5SPILL10_256 <= Tspr5_2_V_1;
                       end 
                      
                  13'sd2357/*2357:xpc10*/:  begin 
                       xpc10 <= 13'sd2358/*2358:xpc10*/;
                       Tsp5SPILL10_256 <= Tspr5_2_V_0;
                       end 
                      
                  13'sd2361/*2361:xpc10*/:  begin 
                       xpc10 <= 13'sd2362/*2362:xpc10*/;
                       Tsf0SPILL12_256 <= 32'sd0;
                       end 
                      
                  13'sd2365/*2365:xpc10*/:  begin 
                       xpc10 <= 13'sd2366/*2366:xpc10*/;
                       Tsf0SPILL10_256 <= 32'sd0;
                       end 
                      
                  13'sd2370/*2370:xpc10*/:  begin 
                       xpc10 <= 13'sd2371/*2371:xpc10*/;
                       Tsf1SPILL12_256 <= 64'h_7fff_ffff_ffff_ffff;
                       end 
                      
                  13'sd2378/*2378:xpc10*/:  begin 
                       xpc10 <= 13'sd2379/*2379:xpc10*/;
                       Tsp7_SPILL_256 <= 64'sh1;
                       end 
                      
                  13'sd2382/*2382:xpc10*/:  begin 
                       xpc10 <= 13'sd2383/*2383:xpc10*/;
                       Tsf1SPILL12_256 <= $signed(64'sh_7ff0_0000_0000_0000+(Tsp7_SPILL_256<<32'sd63));
                       end 
                      
                  13'sd2386/*2386:xpc10*/:  begin 
                       xpc10 <= 13'sd2387/*2387:xpc10*/;
                       Tsp7_SPILL_256 <= 64'sh0;
                       end 
                      
                  13'sd2398/*2398:xpc10*/:  begin 
                       xpc10 <= 13'sd2399/*2399:xpc10*/;
                       Tspr10_2_V_0 <= Tsf1SPILL10_256;
                       end 
                      
                  13'sd2399/*2399:xpc10*/:  begin 
                       xpc10 <= 13'sd2400/*2400:xpc10*/;
                       Tspr10_2_V_1 <= Tsi1SPILL10_256;
                       end 
                      endcase
              if ((32'sd4094/*4094:USA56*/==(64'shfff&(Tspr5_2_V_1>>32'sd51))))  begin if ((13'sd2310/*2310:xpc10*/==xpc10))  xpc10 <= 13'sd2311
                      /*2311:xpc10*/;

                       end 
                   else if ((13'sd2310/*2310:xpc10*/==xpc10))  xpc10 <= 13'sd2359/*2359:xpc10*/;
                      
              case (xpc10)
                  13'sd2304/*2304:xpc10*/:  begin 
                       xpc10 <= 13'sd2305/*2305:xpc10*/;
                       Tsf0SPILL10_256 <= rtl_sign_extend3((32'sd0/*0:USA54*/==(32'sd0/*0:USA52*/==(64'sh7_ffff_ffff_ffff&Tspr5_2_V_0
                      ))));

                       end 
                      
                  13'sd2308/*2308:xpc10*/:  begin 
                       xpc10 <= 13'sd2309/*2309:xpc10*/;
                       Tspr5_2_V_2 <= rtl_unsigned_bitextract4(Tsf0SPILL10_256);
                       end 
                      
                  13'sd2309/*2309:xpc10*/:  begin 
                       xpc10 <= 13'sd2310/*2310:xpc10*/;
                       Tspr5_2_V_3 <= (32'sd0<rtl_sign_extend5(54'sd9007199254740992)+(Tspr5_2_V_1<<32'sd1));
                       end 
                      endcase
              if ((32'sd4094/*4094:USA50*/==(64'shfff&(Tspr5_2_V_0>>32'sd51))))  begin if ((13'sd2300/*2300:xpc10*/==xpc10))  xpc10 <= 13'sd2301
                      /*2301:xpc10*/;

                       end 
                   else if ((13'sd2300/*2300:xpc10*/==xpc10))  xpc10 <= 13'sd2363/*2363:xpc10*/;
                      
              case (xpc10)
                  13'sd2162/*2162:xpc10*/:  begin 
                       xpc10 <= 13'sd2163/*2163:xpc10*/;
                       Tsf0SPILL12_256 <= rtl_sign_extend3((32'sd0/*0:USA160*/==(32'sd0/*0:USA158*/==(64'sh7_ffff_ffff_ffff&Tspr7_3_V_1
                      ))));

                       end 
                      
                  13'sd2166/*2166:xpc10*/:  begin 
                       xpc10 <= 13'sd2167/*2167:xpc10*/;
                       Tspr7_3_V_4 <= rtl_unsigned_bitextract4(Tsf0SPILL12_256);
                       end 
                      
                  13'sd2167/*2167:xpc10*/:  begin 
                       xpc10 <= 13'sd2168/*2168:xpc10*/;
                       Tspr7_3_V_0 <= 64'sh8_0000_0000_0000|Tspr7_3_V_0;
                       end 
                      
                  13'sd2168/*2168:xpc10*/:  begin 
                       xpc10 <= 13'sd2169/*2169:xpc10*/;
                       Tspr7_3_V_1 <= 64'sh8_0000_0000_0000|Tspr7_3_V_1;
                       end 
                      
                  13'sd2169/*2169:xpc10*/:  begin 
                      if (Tspr7_3_V_2 || Tspr7_3_V_4)  begin if (Tspr7_3_V_2 || Tspr7_3_V_4)  xpc10 <= 13'sd2170/*2170:xpc10*/;
                               end 
                          if (!Tspr7_3_V_2 && !Tspr7_3_V_4)  xpc10 <= 13'sd2175/*2175:xpc10*/;
                           end 
                      
                  13'sd2177/*2177:xpc10*/: if (Tspr7_3_V_4)  xpc10 <= 13'sd2178/*2178:xpc10*/;
                       else  xpc10 <= 13'sd2187/*2187:xpc10*/;

                  13'sd2181/*2181:xpc10*/:  begin 
                       xpc10 <= 13'sd2182/*2182:xpc10*/;
                       Tsp7SPILL10_256 <= Tspr7_3_V_1;
                       end 
                      
                  13'sd2185/*2185:xpc10*/:  begin 
                       xpc10 <= 13'sd2186/*2186:xpc10*/;
                       Tss2_SPILL_256 <= Tsp7SPILL10_256;
                       end 
                      
                  13'sd2189/*2189:xpc10*/: if (Tspr7_3_V_2)  xpc10 <= 13'sd2190/*2190:xpc10*/;
                       else  xpc10 <= 13'sd2195/*2195:xpc10*/;

                  13'sd2193/*2193:xpc10*/:  begin 
                       xpc10 <= 13'sd2194/*2194:xpc10*/;
                       Tsp7SPILL10_256 <= Tspr7_3_V_0;
                       end 
                      
                  13'sd2197/*2197:xpc10*/: if (Tspr7_3_V_3)  xpc10 <= 13'sd2198/*2198:xpc10*/;
                       else  xpc10 <= 13'sd2203/*2203:xpc10*/;

                  13'sd2201/*2201:xpc10*/:  begin 
                       xpc10 <= 13'sd2202/*2202:xpc10*/;
                       Tsp7SPILL10_256 <= Tspr7_3_V_1;
                       end 
                      
                  13'sd2205/*2205:xpc10*/:  begin 
                       xpc10 <= 13'sd2206/*2206:xpc10*/;
                       Tsp7SPILL10_256 <= Tspr7_3_V_0;
                       end 
                      
                  13'sd2209/*2209:xpc10*/:  begin 
                       xpc10 <= 13'sd2210/*2210:xpc10*/;
                       Tsf0SPILL12_256 <= 32'sd0;
                       end 
                      
                  13'sd2213/*2213:xpc10*/:  begin 
                       xpc10 <= 13'sd2214/*2214:xpc10*/;
                       Tsf0SPILL10_256 <= 32'sd0;
                       end 
                      
                  13'sd2218/*2218:xpc10*/:  begin 
                       xpc10 <= 13'sd2219/*2219:xpc10*/;
                       Tss2_SPILL_256 <= 64'h_7fff_ffff_ffff_ffff;
                       end 
                      
                  13'sd2226/*2226:xpc10*/:  begin 
                       xpc10 <= 13'sd2227/*2227:xpc10*/;
                       Tssu2_4_V_1 <= 16'sh1;
                       end 
                      
                  13'sd2227/*2227:xpc10*/:  begin 
                       xpc10 <= 13'sd2228/*2228:xpc10*/;
                       Tssu2_4_V_2 <= 16'sh1;
                       end 
                      
                  13'sd2231/*2231:xpc10*/: if ((Tssu2_4_V_5<Tssu2_4_V_4))  xpc10 <= 13'sd2232/*2232:xpc10*/;
                       else  xpc10 <= 13'sd2236/*2236:xpc10*/;

                  13'sd2238/*2238:xpc10*/: if ((Tssu2_4_V_4<Tssu2_4_V_5))  xpc10 <= 13'sd2239/*2239:xpc10*/;
                       else  xpc10 <= 13'sd2243/*2243:xpc10*/;

                  13'sd2249/*2249:xpc10*/:  begin 
                       xpc10 <= 13'sd2250/*2250:xpc10*/;
                       Tsp15_SPILL_256 <= 64'sh0;
                       end 
                      
                  13'sd2250/*2250:xpc10*/:  begin 
                       xpc10 <= 13'sd2251/*2251:xpc10*/;
                       Tss2_SPILL_256 <= 64'h0;
                       end 
                      
                  13'sd2254/*2254:xpc10*/:  begin 
                       xpc10 <= 13'sd2255/*2255:xpc10*/;
                       Tse0SPILL18_256 <= 32'sd0;
                       end 
                      
                  13'sd2258/*2258:xpc10*/:  begin 
                       xpc10 <= 13'sd2259/*2259:xpc10*/;
                       Tse0SPILL16_256 <= 32'sd0;
                       end 
                      
                  13'sd2262/*2262:xpc10*/: if (Tspr2_2_V_2)  xpc10 <= 13'sd2263/*2263:xpc10*/;
                       else  xpc10 <= 13'sd2268/*2268:xpc10*/;

                  13'sd2266/*2266:xpc10*/:  begin 
                       xpc10 <= 13'sd2267/*2267:xpc10*/;
                       Tsp2_SPILL_256 <= Tspr2_2_V_0;
                       end 
                      
                  13'sd2270/*2270:xpc10*/: if (Tspr2_2_V_3)  xpc10 <= 13'sd2271/*2271:xpc10*/;
                       else  xpc10 <= 13'sd2276/*2276:xpc10*/;

                  13'sd2274/*2274:xpc10*/:  begin 
                       xpc10 <= 13'sd2275/*2275:xpc10*/;
                       Tsp2_SPILL_256 <= Tspr2_2_V_1;
                       end 
                      
                  13'sd2278/*2278:xpc10*/:  begin 
                       xpc10 <= 13'sd2279/*2279:xpc10*/;
                       Tsp2_SPILL_256 <= Tspr2_2_V_0;
                       end 
                      
                  13'sd2282/*2282:xpc10*/:  begin 
                       xpc10 <= 13'sd2283/*2283:xpc10*/;
                       Tsf0SPILL12_256 <= 32'sd0;
                       end 
                      
                  13'sd2286/*2286:xpc10*/:  begin 
                       xpc10 <= 13'sd2287/*2287:xpc10*/;
                       Tsf0SPILL10_256 <= 32'sd0;
                       end 
                      
                  13'sd2298/*2298:xpc10*/:  begin 
                       xpc10 <= 13'sd2299/*2299:xpc10*/;
                       Tspr5_2_V_0 <= Tsf1SPILL10_256;
                       end 
                      
                  13'sd2299/*2299:xpc10*/:  begin 
                       xpc10 <= 13'sd2300/*2300:xpc10*/;
                       Tspr5_2_V_1 <= Tsi1SPILL10_256;
                       end 
                      endcase
              if ((32'sd4094/*4094:USA156*/==(64'shfff&(Tspr7_3_V_1>>32'sd51))))  begin if ((13'sd2158/*2158:xpc10*/==xpc10))  xpc10 <= 13'sd2159
                      /*2159:xpc10*/;

                       end 
                   else if ((13'sd2158/*2158:xpc10*/==xpc10))  xpc10 <= 13'sd2207/*2207:xpc10*/;
                      
              case (xpc10)
                  13'sd2152/*2152:xpc10*/:  begin 
                       xpc10 <= 13'sd2153/*2153:xpc10*/;
                       Tsf0SPILL10_256 <= rtl_sign_extend3((32'sd0/*0:USA154*/==(32'sd0/*0:USA152*/==(64'sh7_ffff_ffff_ffff&Tspr7_3_V_0
                      ))));

                       end 
                      
                  13'sd2156/*2156:xpc10*/:  begin 
                       xpc10 <= 13'sd2157/*2157:xpc10*/;
                       Tspr7_3_V_2 <= rtl_unsigned_bitextract4(Tsf0SPILL10_256);
                       end 
                      
                  13'sd2157/*2157:xpc10*/:  begin 
                       xpc10 <= 13'sd2158/*2158:xpc10*/;
                       Tspr7_3_V_3 <= (32'sd0<rtl_sign_extend5(54'sd9007199254740992)+(Tspr7_3_V_1<<32'sd1));
                       end 
                      endcase
              if ((32'sd4094/*4094:USA150*/==(64'shfff&(Tspr7_3_V_0>>32'sd51))))  begin if ((13'sd2148/*2148:xpc10*/==xpc10))  xpc10 <= 13'sd2149
                      /*2149:xpc10*/;

                       end 
                   else if ((13'sd2148/*2148:xpc10*/==xpc10))  xpc10 <= 13'sd2211/*2211:xpc10*/;
                      
              case (xpc10)
                  13'sd2100/*2100:xpc10*/:  begin 
                       xpc10 <= 13'sd2101/*2101:xpc10*/;
                       Tss23_SPILL_258 <= 64'sh1;
                       end 
                      
                  13'sd2101/*2101:xpc10*/:  begin 
                       xpc10 <= 13'sd2102/*2102:xpc10*/;
                       Tss23_SPILL_257 <= Tss23_SPILL_256;
                       end 
                      
                  13'sd2105/*2105:xpc10*/:  begin 
                       xpc10 <= 13'sd2106/*2106:xpc10*/;
                       Tssh23_6_V_0 <= Tss23_SPILL_258|Tss23_SPILL_257;
                       end 
                      
                  13'sd2109/*2109:xpc10*/:  begin 
                       xpc10 <= 13'sd2110/*2110:xpc10*/;
                       Tss23_SPILL_258 <= 64'sh0;
                       end 
                      
                  13'sd2110/*2110:xpc10*/:  begin 
                       xpc10 <= 13'sd2111/*2111:xpc10*/;
                       Tss23_SPILL_257 <= Tss23_SPILL_259;
                       end 
                      
                  13'sd2118/*2118:xpc10*/:  begin 
                       xpc10 <= 13'sd2119/*2119:xpc10*/;
                       Tss23_SPILL_260 <= 64'sh1;
                       end 
                      
                  13'sd2122/*2122:xpc10*/:  begin 
                       xpc10 <= 13'sd2123/*2123:xpc10*/;
                       Tssh23_6_V_0 <= Tss23_SPILL_260;
                       end 
                      
                  13'sd2126/*2126:xpc10*/:  begin 
                       xpc10 <= 13'sd2127/*2127:xpc10*/;
                       Tss23_SPILL_260 <= 64'sh0;
                       end 
                      
                  13'sd2130/*2130:xpc10*/:  begin 
                       xpc10 <= 13'sd2131/*2131:xpc10*/;
                       Tssu2_4_V_4 <= 64'sh_4000_0000_0000_0000|Tssu2_4_V_4;
                       end 
                      
                  13'sd2146/*2146:xpc10*/:  begin 
                       xpc10 <= 13'sd2147/*2147:xpc10*/;
                       Tspr7_3_V_0 <= Tdsi1_5_V_0;
                       end 
                      
                  13'sd2147/*2147:xpc10*/:  begin 
                       xpc10 <= 13'sd2148/*2148:xpc10*/;
                       Tspr7_3_V_1 <= Tdsi1_5_V_1;
                       end 
                      endcase
              if ((32'sd0/*0:USA148*/==(Tssu2_4_V_4<<(32'sd63&rtl_signed_bitextract0(Tssu2_4_V_7)))))  begin if ((13'sd2096/*2096:xpc10*/==
                  xpc10))  xpc10 <= 13'sd2107/*2107:xpc10*/;
                       end 
                   else if ((13'sd2096/*2096:xpc10*/==xpc10))  xpc10 <= 13'sd2097/*2097:xpc10*/;
                      
              case (xpc10)
                  13'sd2050/*2050:xpc10*/:  begin 
                       xpc10 <= 13'sd2051/*2051:xpc10*/;
                       Tsp19_SPILL_256 <= 64'sh1;
                       end 
                      
                  13'sd2054/*2054:xpc10*/:  begin 
                       xpc10 <= 13'sd2055/*2055:xpc10*/;
                       Tss2_SPILL_256 <= $signed(64'sh_7ff0_0000_0000_0000+(Tsp19_SPILL_256<<32'sd63));
                       end 
                      
                  13'sd2058/*2058:xpc10*/:  begin 
                       xpc10 <= 13'sd2059/*2059:xpc10*/;
                       Tsp19_SPILL_256 <= 64'sh0;
                       end 
                      
                  13'sd2066/*2066:xpc10*/:  begin 
                       xpc10 <= 13'sd2067/*2067:xpc10*/;
                       Tssu2_4_V_7 <= 32'sd1+Tssu2_4_V_7;
                       end 
                      
                  13'sd2070/*2070:xpc10*/: if (!(!rtl_signed_bitextract0((0-Tssu2_4_V_7))))  xpc10 <= 13'sd2087/*2087:xpc10*/;
                       else  xpc10 <= 13'sd2071/*2071:xpc10*/;

                  13'sd2074/*2074:xpc10*/:  begin 
                       xpc10 <= 13'sd2075/*2075:xpc10*/;
                       Tssh23_6_V_0 <= Tssu2_4_V_4;
                       end 
                      
                  13'sd2078/*2078:xpc10*/:  begin 
                       xpc10 <= 13'sd2079/*2079:xpc10*/;
                       Tssu2_4_V_4 <= Tssh23_6_V_0;
                       end 
                      
                  13'sd2079/*2079:xpc10*/:  begin 
                       xpc10 <= 13'sd2080/*2080:xpc10*/;
                       Tssu2_4_V_5 <= 64'sh_4000_0000_0000_0000|Tssu2_4_V_5;
                       end 
                      
                  13'sd2083/*2083:xpc10*/:  begin 
                       xpc10 <= 13'sd2084/*2084:xpc10*/;
                       Tssu2_4_V_6 <= Tssu2_4_V_5+(0-Tssu2_4_V_4);
                       end 
                      
                  13'sd2084/*2084:xpc10*/:  begin 
                       xpc10 <= 13'sd2085/*2085:xpc10*/;
                       Tssu2_4_V_3 <= rtl_signed_bitextract0(Tssu2_4_V_2);
                       end 
                      
                  13'sd2085/*2085:xpc10*/:  begin 
                       xpc10 <= 13'sd2086/*2086:xpc10*/;
                       Tssu2_4_V_0 <= (Tssu2_4_V_0==32'sd0/*0:Tssu2.4_V_0*/);
                       end 
                      
                  13'sd2089/*2089:xpc10*/: if ((rtl_signed_bitextract0((0-Tssu2_4_V_7))<32'sd64))  xpc10 <= 13'sd2090/*2090:xpc10*/;
                       else  xpc10 <= 13'sd2112/*2112:xpc10*/;

                  13'sd2093/*2093:xpc10*/:  begin 
                       xpc10 <= 13'sd2094/*2094:xpc10*/;
                       fastspilldup80 <= (Tssu2_4_V_4>>(32'sd63&rtl_signed_bitextract0((0-Tssu2_4_V_7))));
                       end 
                      
                  13'sd2094/*2094:xpc10*/:  begin 
                       xpc10 <= 13'sd2095/*2095:xpc10*/;
                       Tss23_SPILL_259 <= fastspilldup80;
                       end 
                      
                  13'sd2095/*2095:xpc10*/:  begin 
                       xpc10 <= 13'sd2096/*2096:xpc10*/;
                       Tss23_SPILL_256 <= fastspilldup80;
                       end 
                      endcase
              if ((Tssu2_4_V_0==32'sd0/*0:Tssu2.4_V_0*/))  begin if ((13'sd2046/*2046:xpc10*/==xpc10))  xpc10 <= 13'sd2047/*2047:xpc10*/;
                       end 
                   else if ((13'sd2046/*2046:xpc10*/==xpc10))  xpc10 <= 13'sd2056/*2056:xpc10*/;
                      
              case (xpc10)
                  13'sd1991/*1991:xpc10*/:  begin 
                       xpc10 <= 13'sd1992/*1992:xpc10*/;
                       Tsf0SPILL12_256 <= rtl_sign_extend3((32'sd0/*0:USA146*/==(32'sd0/*0:USA144*/==(64'sh7_ffff_ffff_ffff&Tspr18_2_V_1
                      ))));

                       end 
                      
                  13'sd1995/*1995:xpc10*/:  begin 
                       xpc10 <= 13'sd1996/*1996:xpc10*/;
                       Tspr18_2_V_4 <= rtl_unsigned_bitextract4(Tsf0SPILL12_256);
                       end 
                      
                  13'sd1996/*1996:xpc10*/:  begin 
                       xpc10 <= 13'sd1997/*1997:xpc10*/;
                       Tspr18_2_V_0 <= 64'sh8_0000_0000_0000|Tspr18_2_V_0;
                       end 
                      
                  13'sd1997/*1997:xpc10*/:  begin 
                       xpc10 <= 13'sd1998/*1998:xpc10*/;
                       Tspr18_2_V_1 <= 64'sh8_0000_0000_0000|Tspr18_2_V_1;
                       end 
                      
                  13'sd1998/*1998:xpc10*/:  begin 
                      if (Tspr18_2_V_2 || Tspr18_2_V_4)  begin if (Tspr18_2_V_2 || Tspr18_2_V_4)  xpc10 <= 13'sd1999/*1999:xpc10*/;
                               end 
                          if (!Tspr18_2_V_2 && !Tspr18_2_V_4)  xpc10 <= 13'sd2004/*2004:xpc10*/;
                           end 
                      
                  13'sd2006/*2006:xpc10*/: if (Tspr18_2_V_4)  xpc10 <= 13'sd2007/*2007:xpc10*/;
                       else  xpc10 <= 13'sd2016/*2016:xpc10*/;

                  13'sd2010/*2010:xpc10*/:  begin 
                       xpc10 <= 13'sd2011/*2011:xpc10*/;
                       Tsp18SPILL10_256 <= Tspr18_2_V_1;
                       end 
                      
                  13'sd2014/*2014:xpc10*/:  begin 
                       xpc10 <= 13'sd2015/*2015:xpc10*/;
                       Tss2_SPILL_256 <= Tsp18SPILL10_256;
                       end 
                      
                  13'sd2018/*2018:xpc10*/: if (Tspr18_2_V_2)  xpc10 <= 13'sd2019/*2019:xpc10*/;
                       else  xpc10 <= 13'sd2024/*2024:xpc10*/;

                  13'sd2022/*2022:xpc10*/:  begin 
                       xpc10 <= 13'sd2023/*2023:xpc10*/;
                       Tsp18SPILL10_256 <= Tspr18_2_V_0;
                       end 
                      
                  13'sd2026/*2026:xpc10*/: if (Tspr18_2_V_3)  xpc10 <= 13'sd2027/*2027:xpc10*/;
                       else  xpc10 <= 13'sd2032/*2032:xpc10*/;

                  13'sd2030/*2030:xpc10*/:  begin 
                       xpc10 <= 13'sd2031/*2031:xpc10*/;
                       Tsp18SPILL10_256 <= Tspr18_2_V_1;
                       end 
                      
                  13'sd2034/*2034:xpc10*/:  begin 
                       xpc10 <= 13'sd2035/*2035:xpc10*/;
                       Tsp18SPILL10_256 <= Tspr18_2_V_0;
                       end 
                      
                  13'sd2038/*2038:xpc10*/:  begin 
                       xpc10 <= 13'sd2039/*2039:xpc10*/;
                       Tsf0SPILL12_256 <= 32'sd0;
                       end 
                      
                  13'sd2042/*2042:xpc10*/:  begin 
                       xpc10 <= 13'sd2043/*2043:xpc10*/;
                       Tsf0SPILL10_256 <= 32'sd0;
                       end 
                      endcase
              if ((32'sd4094/*4094:USA142*/==(64'shfff&(Tspr18_2_V_1>>32'sd51))))  begin if ((13'sd1987/*1987:xpc10*/==xpc10))  xpc10
                       <= 13'sd1988/*1988:xpc10*/;

                       end 
                   else if ((13'sd1987/*1987:xpc10*/==xpc10))  xpc10 <= 13'sd2036/*2036:xpc10*/;
                      
              case (xpc10)
                  13'sd1981/*1981:xpc10*/:  begin 
                       xpc10 <= 13'sd1982/*1982:xpc10*/;
                       Tsf0SPILL10_256 <= rtl_sign_extend3((32'sd0/*0:USA140*/==(32'sd0/*0:USA138*/==(64'sh7_ffff_ffff_ffff&Tspr18_2_V_0
                      ))));

                       end 
                      
                  13'sd1985/*1985:xpc10*/:  begin 
                       xpc10 <= 13'sd1986/*1986:xpc10*/;
                       Tspr18_2_V_2 <= rtl_unsigned_bitextract4(Tsf0SPILL10_256);
                       end 
                      
                  13'sd1986/*1986:xpc10*/:  begin 
                       xpc10 <= 13'sd1987/*1987:xpc10*/;
                       Tspr18_2_V_3 <= (32'sd0<rtl_sign_extend5(54'sd9007199254740992)+(Tspr18_2_V_1<<32'sd1));
                       end 
                      endcase
              if ((32'sd4094/*4094:USA136*/==(64'shfff&(Tspr18_2_V_0>>32'sd51))))  begin if ((13'sd1977/*1977:xpc10*/==xpc10))  xpc10
                       <= 13'sd1978/*1978:xpc10*/;

                       end 
                   else if ((13'sd1977/*1977:xpc10*/==xpc10))  xpc10 <= 13'sd2040/*2040:xpc10*/;
                      
              case (xpc10)
                  13'sd1975/*1975:xpc10*/:  begin 
                       xpc10 <= 13'sd1976/*1976:xpc10*/;
                       Tspr18_2_V_0 <= Tdsi1_5_V_0;
                       end 
                      
                  13'sd1976/*1976:xpc10*/:  begin 
                       xpc10 <= 13'sd1977/*1977:xpc10*/;
                       Tspr18_2_V_1 <= Tdsi1_5_V_1;
                       end 
                      endcase
              if ((Tssu2_4_V_2==32'sd2047/*2047:Tssu2.4_V_2*/))  begin if ((13'sd1967/*1967:xpc10*/==xpc10))  xpc10 <= 13'sd1968/*1968:xpc10*/;
                       end 
                   else if ((13'sd1967/*1967:xpc10*/==xpc10))  xpc10 <= 13'sd2060/*2060:xpc10*/;
                      
              case (xpc10)
                  13'sd1926/*1926:xpc10*/:  begin 
                       xpc10 <= 13'sd1927/*1927:xpc10*/;
                       Tss32_SPILL_258 <= 64'sh1;
                       end 
                      
                  13'sd1927/*1927:xpc10*/:  begin 
                       xpc10 <= 13'sd1928/*1928:xpc10*/;
                       Tss32_SPILL_257 <= Tss32_SPILL_256;
                       end 
                      
                  13'sd1931/*1931:xpc10*/:  begin 
                       xpc10 <= 13'sd1932/*1932:xpc10*/;
                       Tssh32_5_V_0 <= Tss32_SPILL_258|Tss32_SPILL_257;
                       end 
                      
                  13'sd1935/*1935:xpc10*/:  begin 
                       xpc10 <= 13'sd1936/*1936:xpc10*/;
                       Tss32_SPILL_258 <= 64'sh0;
                       end 
                      
                  13'sd1936/*1936:xpc10*/:  begin 
                       xpc10 <= 13'sd1937/*1937:xpc10*/;
                       Tss32_SPILL_257 <= Tss32_SPILL_259;
                       end 
                      
                  13'sd1944/*1944:xpc10*/:  begin 
                       xpc10 <= 13'sd1945/*1945:xpc10*/;
                       Tss32_SPILL_260 <= 64'sh1;
                       end 
                      
                  13'sd1948/*1948:xpc10*/:  begin 
                       xpc10 <= 13'sd1949/*1949:xpc10*/;
                       Tssh32_5_V_0 <= Tss32_SPILL_260;
                       end 
                      
                  13'sd1952/*1952:xpc10*/:  begin 
                       xpc10 <= 13'sd1953/*1953:xpc10*/;
                       Tss32_SPILL_260 <= 64'sh0;
                       end 
                      
                  13'sd1956/*1956:xpc10*/:  begin 
                       xpc10 <= 13'sd1957/*1957:xpc10*/;
                       Tssu2_4_V_5 <= 64'sh_4000_0000_0000_0000|Tssu2_4_V_5;
                       end 
                      
                  13'sd1960/*1960:xpc10*/: if ((Tssu2_4_V_7<32'sd0))  xpc10 <= 13'sd1961/*1961:xpc10*/;
                       else  xpc10 <= 13'sd2132/*2132:xpc10*/;
              endcase
              if ((32'sd0/*0:USA134*/==(Tssu2_4_V_5<<(32'sd63&rtl_signed_bitextract0((0-Tssu2_4_V_7))))))  begin if ((13'sd1922/*1922:xpc10*/==
                  xpc10))  xpc10 <= 13'sd1933/*1933:xpc10*/;
                       end 
                   else if ((13'sd1922/*1922:xpc10*/==xpc10))  xpc10 <= 13'sd1923/*1923:xpc10*/;
                      
              case (xpc10)
                  13'sd1881/*1881:xpc10*/:  begin 
                       xpc10 <= 13'sd1882/*1882:xpc10*/;
                       Tss18_SPILL_258 <= 64'sh1;
                       end 
                      
                  13'sd1882/*1882:xpc10*/:  begin 
                       xpc10 <= 13'sd1883/*1883:xpc10*/;
                       Tss18_SPILL_257 <= Tss18_SPILL_256;
                       end 
                      
                  13'sd1886/*1886:xpc10*/:  begin 
                       xpc10 <= 13'sd1887/*1887:xpc10*/;
                       Tssh18_7_V_0 <= Tss18_SPILL_258|Tss18_SPILL_257;
                       end 
                      
                  13'sd1890/*1890:xpc10*/:  begin 
                       xpc10 <= 13'sd1891/*1891:xpc10*/;
                       Tss18_SPILL_258 <= 64'sh0;
                       end 
                      
                  13'sd1891/*1891:xpc10*/:  begin 
                       xpc10 <= 13'sd1892/*1892:xpc10*/;
                       Tss18_SPILL_257 <= Tss18_SPILL_259;
                       end 
                      
                  13'sd1899/*1899:xpc10*/:  begin 
                       xpc10 <= 13'sd1900/*1900:xpc10*/;
                       Tss18_SPILL_260 <= 64'sh1;
                       end 
                      
                  13'sd1903/*1903:xpc10*/:  begin 
                       xpc10 <= 13'sd1904/*1904:xpc10*/;
                       Tssh18_7_V_0 <= Tss18_SPILL_260;
                       end 
                      
                  13'sd1907/*1907:xpc10*/:  begin 
                       xpc10 <= 13'sd1908/*1908:xpc10*/;
                       Tss18_SPILL_260 <= 64'sh0;
                       end 
                      
                  13'sd1911/*1911:xpc10*/:  begin 
                       xpc10 <= 13'sd1912/*1912:xpc10*/;
                       Tsco0_2_V_0 <= (Tsco0_2_V_0>>32'sd32);
                       end 
                      
                  13'sd1915/*1915:xpc10*/: if ((rtl_signed_bitextract0(Tssu2_4_V_7)<32'sd64))  xpc10 <= 13'sd1916/*1916:xpc10*/;
                       else  xpc10 <= 13'sd1938/*1938:xpc10*/;

                  13'sd1919/*1919:xpc10*/:  begin 
                       xpc10 <= 13'sd1920/*1920:xpc10*/;
                       fastspilldup82 <= (Tssu2_4_V_5>>(32'sd63&rtl_signed_bitextract0(Tssu2_4_V_7)));
                       end 
                      
                  13'sd1920/*1920:xpc10*/:  begin 
                       xpc10 <= 13'sd1921/*1921:xpc10*/;
                       Tss32_SPILL_259 <= fastspilldup82;
                       end 
                      
                  13'sd1921/*1921:xpc10*/:  begin 
                       xpc10 <= 13'sd1922/*1922:xpc10*/;
                       Tss32_SPILL_256 <= fastspilldup82;
                       end 
                      endcase
              if ((32'sd0/*0:USA162*/==(Tsro0_16_V_1<<(32'sd63&rtl_signed_bitextract0(Tsro0_16_V_0)))))  begin if ((13'sd1877/*1877:xpc10*/==
                  xpc10))  xpc10 <= 13'sd1888/*1888:xpc10*/;
                       end 
                   else if ((13'sd1877/*1877:xpc10*/==xpc10))  xpc10 <= 13'sd1878/*1878:xpc10*/;
                      
              case (xpc10)
                  13'sd1760/*1760:xpc10*/: if ((Tsro0_16_V_1+rtl_sign_extend1(Tsro0_16_V_5)<64'sh0))  xpc10 <= 13'sd1761/*1761:xpc10*/;
                       else  xpc10 <= 13'sd1800/*1800:xpc10*/;

                  13'sd1769/*1769:xpc10*/:  begin 
                       xpc10 <= 13'sd1770/*1770:xpc10*/;
                       Tsp13_SPILL_256 <= 64'sh1;
                       end 
                      
                  13'sd1773/*1773:xpc10*/:  begin 
                       xpc10 <= 13'sd1774/*1774:xpc10*/;
                       fastspilldup84 <= $signed(64'sh_7ff0_0000_0000_0000+(Tsp13_SPILL_256<<32'sd63));
                       end 
                      
                  13'sd1774/*1774:xpc10*/:  begin 
                       xpc10 <= 13'sd1775/*1775:xpc10*/;
                       Tsr0_SPILL_260 <= fastspilldup84;
                       end 
                      
                  13'sd1775/*1775:xpc10*/:  begin 
                       xpc10 <= 13'sd1776/*1776:xpc10*/;
                       Tsr0_SPILL_256 <= fastspilldup84;
                       end 
                      
                  13'sd1776/*1776:xpc10*/: if (!(!Tsro0_16_V_5))  xpc10 <= 13'sd1791/*1791:xpc10*/;
                       else  xpc10 <= 13'sd1777/*1777:xpc10*/;

                  13'sd1780/*1780:xpc10*/:  begin 
                       xpc10 <= 13'sd1781/*1781:xpc10*/;
                       Tsr0_SPILL_258 <= 64'sh1;
                       end 
                      
                  13'sd1781/*1781:xpc10*/:  begin 
                       xpc10 <= 13'sd1782/*1782:xpc10*/;
                       Tsr0_SPILL_257 <= Tsr0_SPILL_256;
                       end 
                      
                  13'sd1785/*1785:xpc10*/:  begin 
                       xpc10 <= 13'sd1786/*1786:xpc10*/;
                       Tsr0_SPILL_259 <= Tsr0_SPILL_257+(0-Tsr0_SPILL_258);
                       end 
                      
                  13'sd1789/*1789:xpc10*/:  begin 
                       xpc10 <= 13'sd1790/*1790:xpc10*/;
                       Tss2_SPILL_256 <= Tsr0_SPILL_259;
                       end 
                      
                  13'sd1793/*1793:xpc10*/:  begin 
                       xpc10 <= 13'sd1794/*1794:xpc10*/;
                       Tsr0_SPILL_258 <= 64'sh0;
                       end 
                      
                  13'sd1794/*1794:xpc10*/:  begin 
                       xpc10 <= 13'sd1795/*1795:xpc10*/;
                       Tsr0_SPILL_257 <= Tsr0_SPILL_260;
                       end 
                      
                  13'sd1798/*1798:xpc10*/:  begin 
                       xpc10 <= 13'sd1799/*1799:xpc10*/;
                       Tsp13_SPILL_256 <= 64'sh0;
                       end 
                      
                  13'sd1802/*1802:xpc10*/: if ((Tsro0_16_V_0<32'sd0))  xpc10 <= 13'sd1803/*1803:xpc10*/;
                       else  xpc10 <= 13'sd1827/*1827:xpc10*/;

                  13'sd1807/*1807:xpc10*/: if (!(!rtl_signed_bitextract0((0-Tsro0_16_V_0))))  xpc10 <= 13'sd1868/*1868:xpc10*/;
                       else  xpc10 <= 13'sd1808/*1808:xpc10*/;

                  13'sd1811/*1811:xpc10*/:  begin 
                       xpc10 <= 13'sd1812/*1812:xpc10*/;
                       Tssh18_7_V_0 <= Tsro0_16_V_1;
                       end 
                      
                  13'sd1815/*1815:xpc10*/:  begin 
                       xpc10 <= 13'sd1816/*1816:xpc10*/;
                       Tsro0_16_V_1 <= Tssh18_7_V_0;
                       end 
                      
                  13'sd1816/*1816:xpc10*/:  begin 
                       xpc10 <= 13'sd1817/*1817:xpc10*/;
                       Tsro0_16_V_0 <= 16'sh0;
                       end 
                      
                  13'sd1817/*1817:xpc10*/:  begin 
                       xpc10 <= 13'sd1818/*1818:xpc10*/;
                       Tsro0_16_V_6 <= rtl_signed_bitextract2(64'sh3ff&Tsro0_16_V_1);
                       end 
                      
                  13'sd1837/*1837:xpc10*/:  begin 
                       xpc10 <= 13'sd1838/*1838:xpc10*/;
                       Tsro0_16_V_1 <= (Tsro0_16_V_1+rtl_sign_extend1(Tsro0_16_V_5)>>32'sd10);
                       end 
                      
                  13'sd1838/*1838:xpc10*/: if (32'sd1&(32'sd0/*0:USA164*/==(32'sd512^Tsro0_16_V_6)))  xpc10 <= 13'sd1839/*1839:xpc10*/;
                       else  xpc10 <= 13'sd1844/*1844:xpc10*/;

                  13'sd1842/*1842:xpc10*/:  begin 
                       xpc10 <= 13'sd1843/*1843:xpc10*/;
                       Tsro0_16_V_1 <= -64'sh2&Tsro0_16_V_1;
                       end 
                      
                  13'sd1850/*1850:xpc10*/:  begin 
                       xpc10 <= 13'sd1851/*1851:xpc10*/;
                       Tsro0_16_V_0 <= 16'sh0;
                       end 
                      
                  13'sd1858/*1858:xpc10*/:  begin 
                       xpc10 <= 13'sd1859/*1859:xpc10*/;
                       Tsp27_SPILL_256 <= 64'sh1;
                       end 
                      
                  13'sd1862/*1862:xpc10*/:  begin 
                       xpc10 <= 13'sd1863/*1863:xpc10*/;
                       Tsr0_SPILL_259 <= Tsro0_16_V_1+(Tsp27_SPILL_256<<32'sd63)+(rtl_sign_extend1(Tsro0_16_V_0)<<32'sd52);
                       end 
                      
                  13'sd1866/*1866:xpc10*/:  begin 
                       xpc10 <= 13'sd1867/*1867:xpc10*/;
                       Tsp27_SPILL_256 <= 64'sh0;
                       end 
                      
                  13'sd1870/*1870:xpc10*/: if ((rtl_signed_bitextract0((0-Tsro0_16_V_0))<32'sd64))  xpc10 <= 13'sd1871/*1871:xpc10*/;
                       else  xpc10 <= 13'sd1893/*1893:xpc10*/;

                  13'sd1874/*1874:xpc10*/:  begin 
                       xpc10 <= 13'sd1875/*1875:xpc10*/;
                       fastspilldup86 <= (Tsro0_16_V_1>>(32'sd63&rtl_signed_bitextract0((0-Tsro0_16_V_0))));
                       end 
                      
                  13'sd1875/*1875:xpc10*/:  begin 
                       xpc10 <= 13'sd1876/*1876:xpc10*/;
                       Tss18_SPILL_259 <= fastspilldup86;
                       end 
                      
                  13'sd1876/*1876:xpc10*/:  begin 
                       xpc10 <= 13'sd1877/*1877:xpc10*/;
                       Tss18_SPILL_256 <= fastspilldup86;
                       end 
                      endcase
              if ((Tsro0_16_V_0==32'sd2045/*2045:Tsro0.16_V_0*/))  begin if ((13'sd1756/*1756:xpc10*/==xpc10))  xpc10 <= 13'sd1757/*1757:xpc10*/;
                       end 
                   else if ((13'sd1756/*1756:xpc10*/==xpc10))  xpc10 <= 13'sd1800/*1800:xpc10*/;
                      
              case (xpc10)
                  13'sd1616/*1616:xpc10*/:  begin 
                       xpc10 <= 13'sd1617/*1617:xpc10*/;
                       Tsf0SPILL12_256 <= rtl_sign_extend3((32'sd0/*0:USA132*/==(32'sd0/*0:USA130*/==(64'sh7_ffff_ffff_ffff&Tspr27_2_V_1
                      ))));

                       end 
                      
                  13'sd1620/*1620:xpc10*/:  begin 
                       xpc10 <= 13'sd1621/*1621:xpc10*/;
                       Tspr27_2_V_4 <= rtl_unsigned_bitextract4(Tsf0SPILL12_256);
                       end 
                      
                  13'sd1621/*1621:xpc10*/:  begin 
                       xpc10 <= 13'sd1622/*1622:xpc10*/;
                       Tspr27_2_V_0 <= 64'sh8_0000_0000_0000|Tspr27_2_V_0;
                       end 
                      
                  13'sd1622/*1622:xpc10*/:  begin 
                       xpc10 <= 13'sd1623/*1623:xpc10*/;
                       Tspr27_2_V_1 <= 64'sh8_0000_0000_0000|Tspr27_2_V_1;
                       end 
                      
                  13'sd1623/*1623:xpc10*/:  begin 
                      if (Tspr27_2_V_2 || Tspr27_2_V_4)  begin if (Tspr27_2_V_2 || Tspr27_2_V_4)  xpc10 <= 13'sd1624/*1624:xpc10*/;
                               end 
                          if (!Tspr27_2_V_2 && !Tspr27_2_V_4)  xpc10 <= 13'sd1629/*1629:xpc10*/;
                           end 
                      
                  13'sd1631/*1631:xpc10*/: if (Tspr27_2_V_4)  xpc10 <= 13'sd1632/*1632:xpc10*/;
                       else  xpc10 <= 13'sd1645/*1645:xpc10*/;

                  13'sd1635/*1635:xpc10*/:  begin 
                       xpc10 <= 13'sd1636/*1636:xpc10*/;
                       Tsp27SPILL10_256 <= Tspr27_2_V_1;
                       end 
                      
                  13'sd1639/*1639:xpc10*/:  begin 
                       xpc10 <= 13'sd1640/*1640:xpc10*/;
                       Tss2_SPILL_256 <= Tsp27SPILL10_256;
                       end 
                      
                  13'sd1643/*1643:xpc10*/:  begin 
                       xpc10 <= 13'sd1644/*1644:xpc10*/;
                       Tsf1SPILL14_256 <= Tss2_SPILL_256;
                       end 
                      
                  13'sd1647/*1647:xpc10*/: if (Tspr27_2_V_2)  xpc10 <= 13'sd1648/*1648:xpc10*/;
                       else  xpc10 <= 13'sd1653/*1653:xpc10*/;

                  13'sd1651/*1651:xpc10*/:  begin 
                       xpc10 <= 13'sd1652/*1652:xpc10*/;
                       Tsp27SPILL10_256 <= Tspr27_2_V_0;
                       end 
                      
                  13'sd1655/*1655:xpc10*/: if (Tspr27_2_V_3)  xpc10 <= 13'sd1656/*1656:xpc10*/;
                       else  xpc10 <= 13'sd1661/*1661:xpc10*/;

                  13'sd1659/*1659:xpc10*/:  begin 
                       xpc10 <= 13'sd1660/*1660:xpc10*/;
                       Tsp27SPILL10_256 <= Tspr27_2_V_1;
                       end 
                      
                  13'sd1663/*1663:xpc10*/:  begin 
                       xpc10 <= 13'sd1664/*1664:xpc10*/;
                       Tsp27SPILL10_256 <= Tspr27_2_V_0;
                       end 
                      
                  13'sd1667/*1667:xpc10*/:  begin 
                       xpc10 <= 13'sd1668/*1668:xpc10*/;
                       Tsf0SPILL12_256 <= 32'sd0;
                       end 
                      
                  13'sd1671/*1671:xpc10*/:  begin 
                       xpc10 <= 13'sd1672/*1672:xpc10*/;
                       Tsf0SPILL10_256 <= 32'sd0;
                       end 
                      
                  13'sd1675/*1675:xpc10*/:  begin 
                       xpc10 <= 13'sd1676/*1676:xpc10*/;
                       Tss2_SPILL_256 <= Tdsi1_5_V_0;
                       end 
                      
                  13'sd1679/*1679:xpc10*/: if (!(!Tssu2_4_V_2))  xpc10 <= 13'sd1954/*1954:xpc10*/;
                       else  xpc10 <= 13'sd1680/*1680:xpc10*/;

                  13'sd1683/*1683:xpc10*/:  begin 
                       xpc10 <= 13'sd1684/*1684:xpc10*/;
                       Tssu2_4_V_7 <= -32'sd1+Tssu2_4_V_7;
                       end 
                      
                  13'sd1687/*1687:xpc10*/: if (!(!rtl_signed_bitextract0(Tssu2_4_V_7)))  xpc10 <= 13'sd1913/*1913:xpc10*/;
                       else  xpc10 <= 13'sd1688/*1688:xpc10*/;

                  13'sd1691/*1691:xpc10*/:  begin 
                       xpc10 <= 13'sd1692/*1692:xpc10*/;
                       Tssh32_5_V_0 <= Tssu2_4_V_5;
                       end 
                      
                  13'sd1695/*1695:xpc10*/:  begin 
                       xpc10 <= 13'sd1696/*1696:xpc10*/;
                       Tssu2_4_V_5 <= Tssh32_5_V_0;
                       end 
                      
                  13'sd1696/*1696:xpc10*/:  begin 
                       xpc10 <= 13'sd1697/*1697:xpc10*/;
                       Tssu2_4_V_4 <= 64'sh_4000_0000_0000_0000|Tssu2_4_V_4;
                       end 
                      
                  13'sd1700/*1700:xpc10*/:  begin 
                       xpc10 <= 13'sd1701/*1701:xpc10*/;
                       Tssu2_4_V_6 <= Tssu2_4_V_4+(0-Tssu2_4_V_5);
                       end 
                      
                  13'sd1701/*1701:xpc10*/:  begin 
                       xpc10 <= 13'sd1702/*1702:xpc10*/;
                       Tssu2_4_V_3 <= rtl_signed_bitextract0(Tssu2_4_V_1);
                       end 
                      
                  13'sd1705/*1705:xpc10*/:  begin 
                       xpc10 <= 13'sd1706/*1706:xpc10*/;
                       Tssu2_4_V_3 <= rtl_signed_bitextract0(-16'sd1+Tssu2_4_V_3);
                       end 
                      
                  13'sd1706/*1706:xpc10*/:  begin 
                       xpc10 <= 13'sd1707/*1707:xpc10*/;
                       Tsco0_2_V_0 <= Tssu2_4_V_6;
                       end 
                      
                  13'sd1707/*1707:xpc10*/:  begin 
                       xpc10 <= 13'sd1708/*1708:xpc10*/;
                       Tsco0_2_V_1 <= 8'h0;
                       end 
                      
                  13'sd1712/*1712:xpc10*/:  begin 
                       xpc10 <= 13'sd1713/*1713:xpc10*/;
                       Tsco0_2_V_1 <= 8'h20;
                       end 
                      
                  13'sd1716/*1716:xpc10*/:  begin 
                       xpc10 <= 13'sd1717/*1717:xpc10*/;
                       Tsco3_7_V_0 <= rtl_unsigned_bitextract6(64'h_ffff_ffff&Tsco0_2_V_0);
                       end 
                      
                  13'sd1717/*1717:xpc10*/:  begin 
                       xpc10 <= 13'sd1718/*1718:xpc10*/;
                       Tsco3_7_V_1 <= 8'h0;
                       end 
                      
                  13'sd1722/*1722:xpc10*/:  begin 
                       xpc10 <= 13'sd1723/*1723:xpc10*/;
                       Tsco3_7_V_1 <= 8'h10;
                       end 
                      
                  13'sd1723/*1723:xpc10*/:  begin 
                       xpc10 <= 13'sd1724/*1724:xpc10*/;
                       Tsco3_7_V_0 <= (Tsco3_7_V_0<<32'sd16);
                       end 
                      
                  13'sd1731/*1731:xpc10*/:  begin 
                       xpc10 <= 13'sd1732/*1732:xpc10*/;
                       Tsco3_7_V_1 <= rtl_unsigned_bitextract7(8'd8+Tsco3_7_V_1);
                       end 
                      
                  13'sd1732/*1732:xpc10*/:  begin 
                       xpc10 <= 13'sd1733/*1733:xpc10*/;
                       Tsco3_7_V_0 <= (Tsco3_7_V_0<<32'sd8);
                       end 
                      
                  13'sd1736/*1736:xpc10*/:  begin 
                       xpc10 <= 13'sd1737/*1737:xpc10*/;
                       Tsco3_7_V_1 <= rtl_unsigned_bitextract7(Tsco3_7_V_1+A_8_US_CC_SCALbx16_ARA0[$unsigned((Tsco3_7_V_0>>32'sd24))]
                      );

                       end 
                      
                  13'sd1737/*1737:xpc10*/:  begin 
                       xpc10 <= 13'sd1738/*1738:xpc10*/;
                       Tsco0_2_V_1 <= rtl_unsigned_bitextract7(Tsco0_2_V_1+Tsco3_7_V_1);
                       end 
                      
                  13'sd1738/*1738:xpc10*/:  begin 
                       xpc10 <= 13'sd1739/*1739:xpc10*/;
                       Tsno34_9_V_0 <= $unsigned(-32'sd1+rtl_sign_extend8(Tsco0_2_V_1));
                       end 
                      
                  13'sd1739/*1739:xpc10*/:  begin 
                       xpc10 <= 13'sd1740/*1740:xpc10*/;
                       Tsro0_16_V_0 <= rtl_signed_bitextract0(rtl_sign_extend9(Tssu2_4_V_3)+(0-Tsno34_9_V_0));
                       end 
                      
                  13'sd1740/*1740:xpc10*/:  begin 
                       xpc10 <= 13'sd1741/*1741:xpc10*/;
                       Tsro0_16_V_1 <= (Tssu2_4_V_6<<(32'sd63&Tsno34_9_V_0));
                       end 
                      
                  13'sd1743/*1743:xpc10*/:  begin 
                       xpc10 <= 13'sd1744/*1744:xpc10*/;
                       Tsro0_16_V_5 <= 16'sh200;
                       end 
                      
                  13'sd1747/*1747:xpc10*/:  begin 
                       xpc10 <= 13'sd1748/*1748:xpc10*/;
                       Tsro0_16_V_6 <= rtl_signed_bitextract2(64'sh3ff&Tsro0_16_V_1);
                       end 
                      
                  13'sd1748/*1748:xpc10*/: if ((Tsro0_16_V_0<32'sd2045))  xpc10 <= 13'sd1827/*1827:xpc10*/;
                       else  xpc10 <= 13'sd1749/*1749:xpc10*/;

                  13'sd1752/*1752:xpc10*/: if ((32'sd2045<Tsro0_16_V_0))  xpc10 <= 13'sd1762/*1762:xpc10*/;
                       else  xpc10 <= 13'sd1753/*1753:xpc10*/;
              endcase
              if ((32'sd4094/*4094:USA128*/==(64'shfff&(Tspr27_2_V_1>>32'sd51))))  begin if ((13'sd1612/*1612:xpc10*/==xpc10))  xpc10
                       <= 13'sd1613/*1613:xpc10*/;

                       end 
                   else if ((13'sd1612/*1612:xpc10*/==xpc10))  xpc10 <= 13'sd1665/*1665:xpc10*/;
                      
              case (xpc10)
                  13'sd1606/*1606:xpc10*/:  begin 
                       xpc10 <= 13'sd1607/*1607:xpc10*/;
                       Tsf0SPILL10_256 <= rtl_sign_extend3((32'sd0/*0:USA126*/==(32'sd0/*0:USA124*/==(64'sh7_ffff_ffff_ffff&Tspr27_2_V_0
                      ))));

                       end 
                      
                  13'sd1610/*1610:xpc10*/:  begin 
                       xpc10 <= 13'sd1611/*1611:xpc10*/;
                       Tspr27_2_V_2 <= rtl_unsigned_bitextract4(Tsf0SPILL10_256);
                       end 
                      
                  13'sd1611/*1611:xpc10*/:  begin 
                       xpc10 <= 13'sd1612/*1612:xpc10*/;
                       Tspr27_2_V_3 <= (32'sd0<rtl_sign_extend5(54'sd9007199254740992)+(Tspr27_2_V_1<<32'sd1));
                       end 
                      endcase
              if ((32'sd4094/*4094:USA122*/==(64'shfff&(Tspr27_2_V_0>>32'sd51))))  begin if ((13'sd1602/*1602:xpc10*/==xpc10))  xpc10
                       <= 13'sd1603/*1603:xpc10*/;

                       end 
                   else if ((13'sd1602/*1602:xpc10*/==xpc10))  xpc10 <= 13'sd1669/*1669:xpc10*/;
                      
              case (xpc10)
                  13'sd1493/*1493:xpc10*/:  begin 
                       xpc10 <= 13'sd1494/*1494:xpc10*/;
                       Tsf0SPILL12_256 <= rtl_sign_extend3((32'sd0/*0:USA116*/==(32'sd0/*0:USA114*/==(64'sh7_ffff_ffff_ffff&Tspr21_3_V_1
                      ))));

                       end 
                      
                  13'sd1497/*1497:xpc10*/:  begin 
                       xpc10 <= 13'sd1498/*1498:xpc10*/;
                       Tspr21_3_V_4 <= rtl_unsigned_bitextract4(Tsf0SPILL12_256);
                       end 
                      
                  13'sd1498/*1498:xpc10*/:  begin 
                       xpc10 <= 13'sd1499/*1499:xpc10*/;
                       Tspr21_3_V_0 <= 64'sh8_0000_0000_0000|Tspr21_3_V_0;
                       end 
                      
                  13'sd1499/*1499:xpc10*/:  begin 
                       xpc10 <= 13'sd1500/*1500:xpc10*/;
                       Tspr21_3_V_1 <= 64'sh8_0000_0000_0000|Tspr21_3_V_1;
                       end 
                      
                  13'sd1500/*1500:xpc10*/:  begin 
                      if (Tspr21_3_V_2 || Tspr21_3_V_4)  begin if (Tspr21_3_V_2 || Tspr21_3_V_4)  xpc10 <= 13'sd1501/*1501:xpc10*/;
                               end 
                          if (!Tspr21_3_V_2 && !Tspr21_3_V_4)  xpc10 <= 13'sd1506/*1506:xpc10*/;
                           end 
                      
                  13'sd1508/*1508:xpc10*/: if (Tspr21_3_V_4)  xpc10 <= 13'sd1509/*1509:xpc10*/;
                       else  xpc10 <= 13'sd1518/*1518:xpc10*/;

                  13'sd1512/*1512:xpc10*/:  begin 
                       xpc10 <= 13'sd1513/*1513:xpc10*/;
                       Tsp21SPILL10_256 <= Tspr21_3_V_1;
                       end 
                      
                  13'sd1516/*1516:xpc10*/:  begin 
                       xpc10 <= 13'sd1517/*1517:xpc10*/;
                       Tsa1_SPILL_256 <= Tsp21SPILL10_256;
                       end 
                      
                  13'sd1520/*1520:xpc10*/: if (Tspr21_3_V_2)  xpc10 <= 13'sd1521/*1521:xpc10*/;
                       else  xpc10 <= 13'sd1526/*1526:xpc10*/;

                  13'sd1524/*1524:xpc10*/:  begin 
                       xpc10 <= 13'sd1525/*1525:xpc10*/;
                       Tsp21SPILL10_256 <= Tspr21_3_V_0;
                       end 
                      
                  13'sd1528/*1528:xpc10*/: if (Tspr21_3_V_3)  xpc10 <= 13'sd1529/*1529:xpc10*/;
                       else  xpc10 <= 13'sd1534/*1534:xpc10*/;

                  13'sd1532/*1532:xpc10*/:  begin 
                       xpc10 <= 13'sd1533/*1533:xpc10*/;
                       Tsp21SPILL10_256 <= Tspr21_3_V_1;
                       end 
                      
                  13'sd1536/*1536:xpc10*/:  begin 
                       xpc10 <= 13'sd1537/*1537:xpc10*/;
                       Tsp21SPILL10_256 <= Tspr21_3_V_0;
                       end 
                      
                  13'sd1540/*1540:xpc10*/:  begin 
                       xpc10 <= 13'sd1541/*1541:xpc10*/;
                       Tsf0SPILL12_256 <= 32'sd0;
                       end 
                      
                  13'sd1544/*1544:xpc10*/:  begin 
                       xpc10 <= 13'sd1545/*1545:xpc10*/;
                       Tsf0SPILL10_256 <= 32'sd0;
                       end 
                      
                  13'sd1548/*1548:xpc10*/:  begin 
                       xpc10 <= 13'sd1549/*1549:xpc10*/;
                       Tsa1_SPILL_256 <= Tdsi1_5_V_0;
                       end 
                      
                  13'sd1560/*1560:xpc10*/:  begin 
                       xpc10 <= 13'sd1561/*1561:xpc10*/;
                       Tsp24_SPILL_256 <= 64'sh1;
                       end 
                      
                  13'sd1564/*1564:xpc10*/:  begin 
                       xpc10 <= 13'sd1565/*1565:xpc10*/;
                       Tsa1_SPILL_256 <= (Tsp24_SPILL_256<<32'sd63)+(Tsad1_3_V_3+Tsad1_3_V_4>>32'sd9);
                       end 
                      
                  13'sd1568/*1568:xpc10*/:  begin 
                       xpc10 <= 13'sd1569/*1569:xpc10*/;
                       Tsp24_SPILL_256 <= 64'sh0;
                       end 
                      
                  13'sd1572/*1572:xpc10*/:  begin 
                       xpc10 <= 13'sd1573/*1573:xpc10*/;
                       Tsad1_3_V_5 <= 64'sh_4000_0000_0000_0000+Tsad1_3_V_3+Tsad1_3_V_4;
                       end 
                      
                  13'sd1573/*1573:xpc10*/:  begin 
                       xpc10 <= 13'sd1574/*1574:xpc10*/;
                       Tsad1_3_V_2 <= rtl_signed_bitextract0(Tsad1_3_V_0);
                       end 
                      
                  13'sd1577/*1577:xpc10*/:  begin 
                       xpc10 <= 13'sd1578/*1578:xpc10*/;
                       Tssu2_4_V_0 <= rtl_unsigned_bitextract12(Tsfl1_39_V_0);
                       end 
                      
                  13'sd1578/*1578:xpc10*/:  begin 
                       xpc10 <= 13'sd1579/*1579:xpc10*/;
                       Tssu2_4_V_4 <= 64'shf_ffff_ffff_ffff&Tdsi1_5_V_0;
                       end 
                      
                  13'sd1579/*1579:xpc10*/:  begin 
                       xpc10 <= 13'sd1580/*1580:xpc10*/;
                       Tssu2_4_V_1 <= rtl_signed_bitextract2(64'sh7ff&(Tdsi1_5_V_0>>32'sd52));
                       end 
                      
                  13'sd1580/*1580:xpc10*/:  begin 
                       xpc10 <= 13'sd1581/*1581:xpc10*/;
                       Tssu2_4_V_5 <= 64'shf_ffff_ffff_ffff&Tdsi1_5_V_1;
                       end 
                      
                  13'sd1581/*1581:xpc10*/:  begin 
                       xpc10 <= 13'sd1582/*1582:xpc10*/;
                       Tssu2_4_V_2 <= rtl_signed_bitextract2(64'sh7ff&(Tdsi1_5_V_1>>32'sd52));
                       end 
                      
                  13'sd1582/*1582:xpc10*/:  begin 
                       xpc10 <= 13'sd1583/*1583:xpc10*/;
                       Tssu2_4_V_7 <= rtl_sign_extend9(Tssu2_4_V_1)+(0-Tssu2_4_V_2);
                       end 
                      
                  13'sd1583/*1583:xpc10*/:  begin 
                       xpc10 <= 13'sd1584/*1584:xpc10*/;
                       Tssu2_4_V_4 <= (Tssu2_4_V_4<<32'sd10);
                       end 
                      
                  13'sd1584/*1584:xpc10*/:  begin 
                       xpc10 <= 13'sd1585/*1585:xpc10*/;
                       Tssu2_4_V_5 <= (Tssu2_4_V_5<<32'sd10);
                       end 
                      
                  13'sd1585/*1585:xpc10*/: if ((32'sd0<Tssu2_4_V_7))  xpc10 <= 13'sd1586/*1586:xpc10*/;
                       else  xpc10 <= 13'sd1958/*1958:xpc10*/;

                  13'sd1600/*1600:xpc10*/:  begin 
                       xpc10 <= 13'sd1601/*1601:xpc10*/;
                       Tspr27_2_V_0 <= Tdsi1_5_V_0;
                       end 
                      
                  13'sd1601/*1601:xpc10*/:  begin 
                       xpc10 <= 13'sd1602/*1602:xpc10*/;
                       Tspr27_2_V_1 <= Tdsi1_5_V_1;
                       end 
                      endcase
              if ((32'sd4094/*4094:USA112*/==(64'shfff&(Tspr21_3_V_1>>32'sd51))))  begin if ((13'sd1489/*1489:xpc10*/==xpc10))  xpc10
                       <= 13'sd1490/*1490:xpc10*/;

                       end 
                   else if ((13'sd1489/*1489:xpc10*/==xpc10))  xpc10 <= 13'sd1538/*1538:xpc10*/;
                      
              case (xpc10)
                  13'sd1483/*1483:xpc10*/:  begin 
                       xpc10 <= 13'sd1484/*1484:xpc10*/;
                       Tsf0SPILL10_256 <= rtl_sign_extend3((32'sd0/*0:USA110*/==(32'sd0/*0:USA108*/==(64'sh7_ffff_ffff_ffff&Tspr21_3_V_0
                      ))));

                       end 
                      
                  13'sd1487/*1487:xpc10*/:  begin 
                       xpc10 <= 13'sd1488/*1488:xpc10*/;
                       Tspr21_3_V_2 <= rtl_unsigned_bitextract4(Tsf0SPILL10_256);
                       end 
                      
                  13'sd1488/*1488:xpc10*/:  begin 
                       xpc10 <= 13'sd1489/*1489:xpc10*/;
                       Tspr21_3_V_3 <= (32'sd0<rtl_sign_extend5(54'sd9007199254740992)+(Tspr21_3_V_1<<32'sd1));
                       end 
                      endcase
              if ((32'sd4094/*4094:USA106*/==(64'shfff&(Tspr21_3_V_0>>32'sd51))))  begin if ((13'sd1479/*1479:xpc10*/==xpc10))  xpc10
                       <= 13'sd1480/*1480:xpc10*/;

                       end 
                   else if ((13'sd1479/*1479:xpc10*/==xpc10))  xpc10 <= 13'sd1542/*1542:xpc10*/;
                      
              case (xpc10)
                  13'sd1431/*1431:xpc10*/:  begin 
                       xpc10 <= 13'sd1432/*1432:xpc10*/;
                       Tss17_SPILL_258 <= 64'sh1;
                       end 
                      
                  13'sd1432/*1432:xpc10*/:  begin 
                       xpc10 <= 13'sd1433/*1433:xpc10*/;
                       Tss17_SPILL_257 <= Tss17_SPILL_256;
                       end 
                      
                  13'sd1436/*1436:xpc10*/:  begin 
                       xpc10 <= 13'sd1437/*1437:xpc10*/;
                       Tssh17_6_V_0 <= Tss17_SPILL_258|Tss17_SPILL_257;
                       end 
                      
                  13'sd1440/*1440:xpc10*/:  begin 
                       xpc10 <= 13'sd1441/*1441:xpc10*/;
                       Tss17_SPILL_258 <= 64'sh0;
                       end 
                      
                  13'sd1441/*1441:xpc10*/:  begin 
                       xpc10 <= 13'sd1442/*1442:xpc10*/;
                       Tss17_SPILL_257 <= Tss17_SPILL_259;
                       end 
                      
                  13'sd1449/*1449:xpc10*/:  begin 
                       xpc10 <= 13'sd1450/*1450:xpc10*/;
                       Tss17_SPILL_260 <= 64'sh1;
                       end 
                      
                  13'sd1453/*1453:xpc10*/:  begin 
                       xpc10 <= 13'sd1454/*1454:xpc10*/;
                       Tssh17_6_V_0 <= Tss17_SPILL_260;
                       end 
                      
                  13'sd1457/*1457:xpc10*/:  begin 
                       xpc10 <= 13'sd1458/*1458:xpc10*/;
                       Tss17_SPILL_260 <= 64'sh0;
                       end 
                      
                  13'sd1461/*1461:xpc10*/:  begin 
                       xpc10 <= 13'sd1462/*1462:xpc10*/;
                       Tsad1_3_V_3 <= 64'sh_2000_0000_0000_0000|Tsad1_3_V_3;
                       end 
                      
                  13'sd1477/*1477:xpc10*/:  begin 
                       xpc10 <= 13'sd1478/*1478:xpc10*/;
                       Tspr21_3_V_0 <= Tdsi1_5_V_0;
                       end 
                      
                  13'sd1478/*1478:xpc10*/:  begin 
                       xpc10 <= 13'sd1479/*1479:xpc10*/;
                       Tspr21_3_V_1 <= Tdsi1_5_V_1;
                       end 
                      endcase
              if ((32'sd0/*0:USA104*/==(Tsad1_3_V_3<<(32'sd63&rtl_signed_bitextract0(Tsad1_3_V_6)))))  begin if ((13'sd1427/*1427:xpc10*/==
                  xpc10))  xpc10 <= 13'sd1438/*1438:xpc10*/;
                       end 
                   else if ((13'sd1427/*1427:xpc10*/==xpc10))  xpc10 <= 13'sd1428/*1428:xpc10*/;
                      
              case (xpc10)
                  13'sd1328/*1328:xpc10*/:  begin 
                       xpc10 <= 13'sd1329/*1329:xpc10*/;
                       Tsf0SPILL12_256 <= rtl_sign_extend3((32'sd0/*0:USA102*/==(32'sd0/*0:USA100*/==(64'sh7_ffff_ffff_ffff&Tspr12_2_V_1
                      ))));

                       end 
                      
                  13'sd1332/*1332:xpc10*/:  begin 
                       xpc10 <= 13'sd1333/*1333:xpc10*/;
                       Tspr12_2_V_4 <= rtl_unsigned_bitextract4(Tsf0SPILL12_256);
                       end 
                      
                  13'sd1333/*1333:xpc10*/:  begin 
                       xpc10 <= 13'sd1334/*1334:xpc10*/;
                       Tspr12_2_V_0 <= 64'sh8_0000_0000_0000|Tspr12_2_V_0;
                       end 
                      
                  13'sd1334/*1334:xpc10*/:  begin 
                       xpc10 <= 13'sd1335/*1335:xpc10*/;
                       Tspr12_2_V_1 <= 64'sh8_0000_0000_0000|Tspr12_2_V_1;
                       end 
                      
                  13'sd1335/*1335:xpc10*/:  begin 
                      if (Tspr12_2_V_2 || Tspr12_2_V_4)  begin if (Tspr12_2_V_2 || Tspr12_2_V_4)  xpc10 <= 13'sd1336/*1336:xpc10*/;
                               end 
                          if (!Tspr12_2_V_2 && !Tspr12_2_V_4)  xpc10 <= 13'sd1341/*1341:xpc10*/;
                           end 
                      
                  13'sd1343/*1343:xpc10*/: if (Tspr12_2_V_4)  xpc10 <= 13'sd1344/*1344:xpc10*/;
                       else  xpc10 <= 13'sd1353/*1353:xpc10*/;

                  13'sd1347/*1347:xpc10*/:  begin 
                       xpc10 <= 13'sd1348/*1348:xpc10*/;
                       Tsp12_SPILL_256 <= Tspr12_2_V_1;
                       end 
                      
                  13'sd1351/*1351:xpc10*/:  begin 
                       xpc10 <= 13'sd1352/*1352:xpc10*/;
                       Tsa1_SPILL_256 <= Tsp12_SPILL_256;
                       end 
                      
                  13'sd1355/*1355:xpc10*/: if (Tspr12_2_V_2)  xpc10 <= 13'sd1356/*1356:xpc10*/;
                       else  xpc10 <= 13'sd1361/*1361:xpc10*/;

                  13'sd1359/*1359:xpc10*/:  begin 
                       xpc10 <= 13'sd1360/*1360:xpc10*/;
                       Tsp12_SPILL_256 <= Tspr12_2_V_0;
                       end 
                      
                  13'sd1363/*1363:xpc10*/: if (Tspr12_2_V_3)  xpc10 <= 13'sd1364/*1364:xpc10*/;
                       else  xpc10 <= 13'sd1369/*1369:xpc10*/;

                  13'sd1367/*1367:xpc10*/:  begin 
                       xpc10 <= 13'sd1368/*1368:xpc10*/;
                       Tsp12_SPILL_256 <= Tspr12_2_V_1;
                       end 
                      
                  13'sd1371/*1371:xpc10*/:  begin 
                       xpc10 <= 13'sd1372/*1372:xpc10*/;
                       Tsp12_SPILL_256 <= Tspr12_2_V_0;
                       end 
                      
                  13'sd1375/*1375:xpc10*/:  begin 
                       xpc10 <= 13'sd1376/*1376:xpc10*/;
                       Tsf0SPILL12_256 <= 32'sd0;
                       end 
                      
                  13'sd1379/*1379:xpc10*/:  begin 
                       xpc10 <= 13'sd1380/*1380:xpc10*/;
                       Tsf0SPILL10_256 <= 32'sd0;
                       end 
                      
                  13'sd1387/*1387:xpc10*/:  begin 
                       xpc10 <= 13'sd1388/*1388:xpc10*/;
                       Tsp13SPILL10_256 <= 64'sh1;
                       end 
                      
                  13'sd1391/*1391:xpc10*/:  begin 
                       xpc10 <= 13'sd1392/*1392:xpc10*/;
                       Tsa1_SPILL_256 <= $signed(64'sh_7ff0_0000_0000_0000+(Tsp13SPILL10_256<<32'sd63));
                       end 
                      
                  13'sd1395/*1395:xpc10*/:  begin 
                       xpc10 <= 13'sd1396/*1396:xpc10*/;
                       Tsp13SPILL10_256 <= 64'sh0;
                       end 
                      
                  13'sd1403/*1403:xpc10*/:  begin 
                       xpc10 <= 13'sd1404/*1404:xpc10*/;
                       Tsad1_3_V_6 <= 32'sd1+Tsad1_3_V_6;
                       end 
                      
                  13'sd1407/*1407:xpc10*/: if (!(!rtl_signed_bitextract0((0-Tsad1_3_V_6))))  xpc10 <= 13'sd1418/*1418:xpc10*/;
                       else  xpc10 <= 13'sd1408/*1408:xpc10*/;

                  13'sd1411/*1411:xpc10*/:  begin 
                       xpc10 <= 13'sd1412/*1412:xpc10*/;
                       Tssh17_6_V_0 <= Tsad1_3_V_3;
                       end 
                      
                  13'sd1415/*1415:xpc10*/:  begin 
                       xpc10 <= 13'sd1416/*1416:xpc10*/;
                       Tsad1_3_V_3 <= Tssh17_6_V_0;
                       end 
                      
                  13'sd1416/*1416:xpc10*/:  begin 
                       xpc10 <= 13'sd1417/*1417:xpc10*/;
                       Tsad1_3_V_2 <= rtl_signed_bitextract0(Tsad1_3_V_1);
                       end 
                      
                  13'sd1420/*1420:xpc10*/: if ((rtl_signed_bitextract0((0-Tsad1_3_V_6))<32'sd64))  xpc10 <= 13'sd1421/*1421:xpc10*/;
                       else  xpc10 <= 13'sd1443/*1443:xpc10*/;

                  13'sd1424/*1424:xpc10*/:  begin 
                       xpc10 <= 13'sd1425/*1425:xpc10*/;
                       fastspilldup74 <= (Tsad1_3_V_3>>(32'sd63&rtl_signed_bitextract0((0-Tsad1_3_V_6))));
                       end 
                      
                  13'sd1425/*1425:xpc10*/:  begin 
                       xpc10 <= 13'sd1426/*1426:xpc10*/;
                       Tss17_SPILL_259 <= fastspilldup74;
                       end 
                      
                  13'sd1426/*1426:xpc10*/:  begin 
                       xpc10 <= 13'sd1427/*1427:xpc10*/;
                       Tss17_SPILL_256 <= fastspilldup74;
                       end 
                      endcase
              if ((32'sd4094/*4094:USA98*/==(64'shfff&(Tspr12_2_V_1>>32'sd51))))  begin if ((13'sd1324/*1324:xpc10*/==xpc10))  xpc10 <= 13'sd1325
                      /*1325:xpc10*/;

                       end 
                   else if ((13'sd1324/*1324:xpc10*/==xpc10))  xpc10 <= 13'sd1373/*1373:xpc10*/;
                      
              case (xpc10)
                  13'sd1318/*1318:xpc10*/:  begin 
                       xpc10 <= 13'sd1319/*1319:xpc10*/;
                       Tsf0SPILL10_256 <= rtl_sign_extend3((32'sd0/*0:USA96*/==(32'sd0/*0:USA94*/==(64'sh7_ffff_ffff_ffff&Tspr12_2_V_0
                      ))));

                       end 
                      
                  13'sd1322/*1322:xpc10*/:  begin 
                       xpc10 <= 13'sd1323/*1323:xpc10*/;
                       Tspr12_2_V_2 <= rtl_unsigned_bitextract4(Tsf0SPILL10_256);
                       end 
                      
                  13'sd1323/*1323:xpc10*/:  begin 
                       xpc10 <= 13'sd1324/*1324:xpc10*/;
                       Tspr12_2_V_3 <= (32'sd0<rtl_sign_extend5(54'sd9007199254740992)+(Tspr12_2_V_1<<32'sd1));
                       end 
                      endcase
              if ((32'sd4094/*4094:USA92*/==(64'shfff&(Tspr12_2_V_0>>32'sd51))))  begin if ((13'sd1314/*1314:xpc10*/==xpc10))  xpc10 <= 13'sd1315
                      /*1315:xpc10*/;

                       end 
                   else if ((13'sd1314/*1314:xpc10*/==xpc10))  xpc10 <= 13'sd1377/*1377:xpc10*/;
                      
              case (xpc10)
                  13'sd1312/*1312:xpc10*/:  begin 
                       xpc10 <= 13'sd1313/*1313:xpc10*/;
                       Tspr12_2_V_0 <= Tdsi1_5_V_0;
                       end 
                      
                  13'sd1313/*1313:xpc10*/:  begin 
                       xpc10 <= 13'sd1314/*1314:xpc10*/;
                       Tspr12_2_V_1 <= Tdsi1_5_V_1;
                       end 
                      endcase
              if ((Tsad1_3_V_1==32'sd2047/*2047:Tsad1.3_V_1*/))  begin if ((13'sd1304/*1304:xpc10*/==xpc10))  xpc10 <= 13'sd1305/*1305:xpc10*/;
                       end 
                   else if ((13'sd1304/*1304:xpc10*/==xpc10))  xpc10 <= 13'sd1397/*1397:xpc10*/;
                      
              case (xpc10)
                  13'sd1266/*1266:xpc10*/:  begin 
                       xpc10 <= 13'sd1267/*1267:xpc10*/;
                       Tss8_SPILL_258 <= 64'sh1;
                       end 
                      
                  13'sd1267/*1267:xpc10*/:  begin 
                       xpc10 <= 13'sd1268/*1268:xpc10*/;
                       Tss8_SPILL_257 <= Tss8_SPILL_256;
                       end 
                      
                  13'sd1271/*1271:xpc10*/:  begin 
                       xpc10 <= 13'sd1272/*1272:xpc10*/;
                       Tssh8_5_V_0 <= Tss8_SPILL_258|Tss8_SPILL_257;
                       end 
                      
                  13'sd1275/*1275:xpc10*/:  begin 
                       xpc10 <= 13'sd1276/*1276:xpc10*/;
                       Tss8_SPILL_258 <= 64'sh0;
                       end 
                      
                  13'sd1276/*1276:xpc10*/:  begin 
                       xpc10 <= 13'sd1277/*1277:xpc10*/;
                       Tss8_SPILL_257 <= Tss8_SPILL_259;
                       end 
                      
                  13'sd1284/*1284:xpc10*/:  begin 
                       xpc10 <= 13'sd1285/*1285:xpc10*/;
                       Tss8_SPILL_260 <= 64'sh1;
                       end 
                      
                  13'sd1288/*1288:xpc10*/:  begin 
                       xpc10 <= 13'sd1289/*1289:xpc10*/;
                       Tssh8_5_V_0 <= Tss8_SPILL_260;
                       end 
                      
                  13'sd1292/*1292:xpc10*/:  begin 
                       xpc10 <= 13'sd1293/*1293:xpc10*/;
                       Tss8_SPILL_260 <= 64'sh0;
                       end 
                      
                  13'sd1296/*1296:xpc10*/:  begin 
                       xpc10 <= 13'sd1297/*1297:xpc10*/;
                       Tsad1_3_V_4 <= 64'sh_2000_0000_0000_0000|Tsad1_3_V_4;
                       end 
                      
                  13'sd1300/*1300:xpc10*/: if ((Tsad1_3_V_6<32'sd0))  xpc10 <= 13'sd1301/*1301:xpc10*/;
                       else  xpc10 <= 13'sd1463/*1463:xpc10*/;
              endcase
              if ((32'sd0/*0:USA90*/==(Tsad1_3_V_4<<(32'sd63&rtl_signed_bitextract0((0-Tsad1_3_V_6))))))  begin if ((13'sd1262/*1262:xpc10*/==
                  xpc10))  xpc10 <= 13'sd1273/*1273:xpc10*/;
                       end 
                   else if ((13'sd1262/*1262:xpc10*/==xpc10))  xpc10 <= 13'sd1263/*1263:xpc10*/;
                      
              case (xpc10)
                  13'sd1225/*1225:xpc10*/:  begin 
                       xpc10 <= 13'sd1226/*1226:xpc10*/;
                       Tss18_SPILL_258 <= 64'sh1;
                       end 
                      
                  13'sd1226/*1226:xpc10*/:  begin 
                       xpc10 <= 13'sd1227/*1227:xpc10*/;
                       Tss18_SPILL_257 <= Tss18_SPILL_256;
                       end 
                      
                  13'sd1230/*1230:xpc10*/:  begin 
                       xpc10 <= 13'sd1231/*1231:xpc10*/;
                       Tssh18_7_V_0 <= Tss18_SPILL_258|Tss18_SPILL_257;
                       end 
                      
                  13'sd1234/*1234:xpc10*/:  begin 
                       xpc10 <= 13'sd1235/*1235:xpc10*/;
                       Tss18_SPILL_258 <= 64'sh0;
                       end 
                      
                  13'sd1235/*1235:xpc10*/:  begin 
                       xpc10 <= 13'sd1236/*1236:xpc10*/;
                       Tss18_SPILL_257 <= Tss18_SPILL_259;
                       end 
                      
                  13'sd1243/*1243:xpc10*/:  begin 
                       xpc10 <= 13'sd1244/*1244:xpc10*/;
                       Tss18_SPILL_260 <= 64'sh1;
                       end 
                      
                  13'sd1247/*1247:xpc10*/:  begin 
                       xpc10 <= 13'sd1248/*1248:xpc10*/;
                       Tssh18_7_V_0 <= Tss18_SPILL_260;
                       end 
                      
                  13'sd1251/*1251:xpc10*/:  begin 
                       xpc10 <= 13'sd1252/*1252:xpc10*/;
                       Tss18_SPILL_260 <= 64'sh0;
                       end 
                      
                  13'sd1255/*1255:xpc10*/: if ((rtl_signed_bitextract0(Tsad1_3_V_6)<32'sd64))  xpc10 <= 13'sd1256/*1256:xpc10*/;
                       else  xpc10 <= 13'sd1278/*1278:xpc10*/;

                  13'sd1259/*1259:xpc10*/:  begin 
                       xpc10 <= 13'sd1260/*1260:xpc10*/;
                       fastspilldup72 <= (Tsad1_3_V_4>>(32'sd63&rtl_signed_bitextract0(Tsad1_3_V_6)));
                       end 
                      
                  13'sd1260/*1260:xpc10*/:  begin 
                       xpc10 <= 13'sd1261/*1261:xpc10*/;
                       Tss8_SPILL_259 <= fastspilldup72;
                       end 
                      
                  13'sd1261/*1261:xpc10*/:  begin 
                       xpc10 <= 13'sd1262/*1262:xpc10*/;
                       Tss8_SPILL_256 <= fastspilldup72;
                       end 
                      endcase
              if ((32'sd0/*0:USA118*/==(Tsro28_4_V_1<<(32'sd63&rtl_signed_bitextract0(Tsro28_4_V_0)))))  begin if ((13'sd1221/*1221:xpc10*/==
                  xpc10))  xpc10 <= 13'sd1232/*1232:xpc10*/;
                       end 
                   else if ((13'sd1221/*1221:xpc10*/==xpc10))  xpc10 <= 13'sd1222/*1222:xpc10*/;
                      
              case (xpc10)
                  13'sd1104/*1104:xpc10*/: if ((Tsro28_4_V_1+rtl_sign_extend1(Tsro28_4_V_5)<64'sh0))  xpc10 <= 13'sd1105/*1105:xpc10*/;
                       else  xpc10 <= 13'sd1144/*1144:xpc10*/;

                  13'sd1113/*1113:xpc10*/:  begin 
                       xpc10 <= 13'sd1114/*1114:xpc10*/;
                       Tsp13_SPILL_256 <= 64'sh1;
                       end 
                      
                  13'sd1117/*1117:xpc10*/:  begin 
                       xpc10 <= 13'sd1118/*1118:xpc10*/;
                       fastspilldup76 <= $signed(64'sh_7ff0_0000_0000_0000+(Tsp13_SPILL_256<<32'sd63));
                       end 
                      
                  13'sd1118/*1118:xpc10*/:  begin 
                       xpc10 <= 13'sd1119/*1119:xpc10*/;
                       Tsr28_SPILL_260 <= fastspilldup76;
                       end 
                      
                  13'sd1119/*1119:xpc10*/:  begin 
                       xpc10 <= 13'sd1120/*1120:xpc10*/;
                       Tsr28_SPILL_256 <= fastspilldup76;
                       end 
                      
                  13'sd1120/*1120:xpc10*/: if (!(!Tsro28_4_V_5))  xpc10 <= 13'sd1135/*1135:xpc10*/;
                       else  xpc10 <= 13'sd1121/*1121:xpc10*/;

                  13'sd1124/*1124:xpc10*/:  begin 
                       xpc10 <= 13'sd1125/*1125:xpc10*/;
                       Tsr28_SPILL_258 <= 64'sh1;
                       end 
                      
                  13'sd1125/*1125:xpc10*/:  begin 
                       xpc10 <= 13'sd1126/*1126:xpc10*/;
                       Tsr28_SPILL_257 <= Tsr28_SPILL_256;
                       end 
                      
                  13'sd1129/*1129:xpc10*/:  begin 
                       xpc10 <= 13'sd1130/*1130:xpc10*/;
                       Tsr28_SPILL_259 <= Tsr28_SPILL_257+(0-Tsr28_SPILL_258);
                       end 
                      
                  13'sd1133/*1133:xpc10*/:  begin 
                       xpc10 <= 13'sd1134/*1134:xpc10*/;
                       Tsa1_SPILL_256 <= Tsr28_SPILL_259;
                       end 
                      
                  13'sd1137/*1137:xpc10*/:  begin 
                       xpc10 <= 13'sd1138/*1138:xpc10*/;
                       Tsr28_SPILL_258 <= 64'sh0;
                       end 
                      
                  13'sd1138/*1138:xpc10*/:  begin 
                       xpc10 <= 13'sd1139/*1139:xpc10*/;
                       Tsr28_SPILL_257 <= Tsr28_SPILL_260;
                       end 
                      
                  13'sd1142/*1142:xpc10*/:  begin 
                       xpc10 <= 13'sd1143/*1143:xpc10*/;
                       Tsp13_SPILL_256 <= 64'sh0;
                       end 
                      
                  13'sd1146/*1146:xpc10*/: if ((Tsro28_4_V_0<32'sd0))  xpc10 <= 13'sd1147/*1147:xpc10*/;
                       else  xpc10 <= 13'sd1171/*1171:xpc10*/;

                  13'sd1151/*1151:xpc10*/: if (!(!rtl_signed_bitextract0((0-Tsro28_4_V_0))))  xpc10 <= 13'sd1212/*1212:xpc10*/;
                       else  xpc10 <= 13'sd1152/*1152:xpc10*/;

                  13'sd1155/*1155:xpc10*/:  begin 
                       xpc10 <= 13'sd1156/*1156:xpc10*/;
                       Tssh18_7_V_0 <= Tsro28_4_V_1;
                       end 
                      
                  13'sd1159/*1159:xpc10*/:  begin 
                       xpc10 <= 13'sd1160/*1160:xpc10*/;
                       Tsro28_4_V_1 <= Tssh18_7_V_0;
                       end 
                      
                  13'sd1160/*1160:xpc10*/:  begin 
                       xpc10 <= 13'sd1161/*1161:xpc10*/;
                       Tsro28_4_V_0 <= 16'sh0;
                       end 
                      
                  13'sd1161/*1161:xpc10*/:  begin 
                       xpc10 <= 13'sd1162/*1162:xpc10*/;
                       Tsro28_4_V_6 <= rtl_signed_bitextract2(64'sh3ff&Tsro28_4_V_1);
                       end 
                      
                  13'sd1181/*1181:xpc10*/:  begin 
                       xpc10 <= 13'sd1182/*1182:xpc10*/;
                       Tsro28_4_V_1 <= (Tsro28_4_V_1+rtl_sign_extend1(Tsro28_4_V_5)>>32'sd10);
                       end 
                      
                  13'sd1182/*1182:xpc10*/: if (32'sd1&(32'sd0/*0:USA120*/==(32'sd512^Tsro28_4_V_6)))  xpc10 <= 13'sd1183/*1183:xpc10*/;
                       else  xpc10 <= 13'sd1188/*1188:xpc10*/;

                  13'sd1186/*1186:xpc10*/:  begin 
                       xpc10 <= 13'sd1187/*1187:xpc10*/;
                       Tsro28_4_V_1 <= -64'sh2&Tsro28_4_V_1;
                       end 
                      
                  13'sd1194/*1194:xpc10*/:  begin 
                       xpc10 <= 13'sd1195/*1195:xpc10*/;
                       Tsro28_4_V_0 <= 16'sh0;
                       end 
                      
                  13'sd1202/*1202:xpc10*/:  begin 
                       xpc10 <= 13'sd1203/*1203:xpc10*/;
                       Tsp27_SPILL_256 <= 64'sh1;
                       end 
                      
                  13'sd1206/*1206:xpc10*/:  begin 
                       xpc10 <= 13'sd1207/*1207:xpc10*/;
                       Tsr28_SPILL_259 <= Tsro28_4_V_1+(Tsp27_SPILL_256<<32'sd63)+(rtl_sign_extend1(Tsro28_4_V_0)<<32'sd52);
                       end 
                      
                  13'sd1210/*1210:xpc10*/:  begin 
                       xpc10 <= 13'sd1211/*1211:xpc10*/;
                       Tsp27_SPILL_256 <= 64'sh0;
                       end 
                      
                  13'sd1214/*1214:xpc10*/: if ((rtl_signed_bitextract0((0-Tsro28_4_V_0))<32'sd64))  xpc10 <= 13'sd1215/*1215:xpc10*/;
                       else  xpc10 <= 13'sd1237/*1237:xpc10*/;

                  13'sd1218/*1218:xpc10*/:  begin 
                       xpc10 <= 13'sd1219/*1219:xpc10*/;
                       fastspilldup78 <= (Tsro28_4_V_1>>(32'sd63&rtl_signed_bitextract0((0-Tsro28_4_V_0))));
                       end 
                      
                  13'sd1219/*1219:xpc10*/:  begin 
                       xpc10 <= 13'sd1220/*1220:xpc10*/;
                       Tss18_SPILL_259 <= fastspilldup78;
                       end 
                      
                  13'sd1220/*1220:xpc10*/:  begin 
                       xpc10 <= 13'sd1221/*1221:xpc10*/;
                       Tss18_SPILL_256 <= fastspilldup78;
                       end 
                      endcase
              if ((Tsro28_4_V_0==32'sd2045/*2045:Tsro28.4_V_0*/))  begin if ((13'sd1100/*1100:xpc10*/==xpc10))  xpc10 <= 13'sd1101/*1101:xpc10*/;
                       end 
                   else if ((13'sd1100/*1100:xpc10*/==xpc10))  xpc10 <= 13'sd1144/*1144:xpc10*/;
                      
              case (xpc10)
                  13'sd1002/*1002:xpc10*/:  begin 
                       xpc10 <= 13'sd1003/*1003:xpc10*/;
                       Tsf0SPILL14_258 <= $unsigned(Tsfl0_3_V_0^(64'sh_3ee4_f8b5_88e3_68f1<(64'sh_7fff_ffff_ffff_ffff&Tdsi1_5_V_1)));
                       end 
                      
                  13'sd1006/*1006:xpc10*/:  begin 
                       xpc10 <= 13'sd1007/*1007:xpc10*/;
                       Tsf0SPILL14_256 <= Tsf0SPILL14_258;
                       end 
                      
                  13'sd1010/*1010:xpc10*/:  begin 
                       xpc10 <= 13'sd1011/*1011:xpc10*/;
                       Tsf0SPILL14_258 <= 32'sd1;
                       end 
                      
                  13'sd1014/*1014:xpc10*/:  begin 
                       xpc10 <= 13'sd1015/*1015:xpc10*/;
                       Tse5SPILL10_256 <= 32'sd0;
                       end 
                      
                  13'sd1018/*1018:xpc10*/: if (Tspr3_2_V_2)  xpc10 <= 13'sd1019/*1019:xpc10*/;
                       else  xpc10 <= 13'sd1024/*1024:xpc10*/;

                  13'sd1022/*1022:xpc10*/:  begin 
                       xpc10 <= 13'sd1023/*1023:xpc10*/;
                       Tsp3_SPILL_256 <= Tspr3_2_V_0;
                       end 
                      
                  13'sd1026/*1026:xpc10*/: if (Tspr3_2_V_3)  xpc10 <= 13'sd1027/*1027:xpc10*/;
                       else  xpc10 <= 13'sd1032/*1032:xpc10*/;

                  13'sd1030/*1030:xpc10*/:  begin 
                       xpc10 <= 13'sd1031/*1031:xpc10*/;
                       Tsp3_SPILL_256 <= Tspr3_2_V_1;
                       end 
                      
                  13'sd1034/*1034:xpc10*/:  begin 
                       xpc10 <= 13'sd1035/*1035:xpc10*/;
                       Tsp3_SPILL_256 <= Tspr3_2_V_0;
                       end 
                      
                  13'sd1038/*1038:xpc10*/:  begin 
                       xpc10 <= 13'sd1039/*1039:xpc10*/;
                       Tsf0SPILL12_256 <= 32'sd0;
                       end 
                      
                  13'sd1042/*1042:xpc10*/:  begin 
                       xpc10 <= 13'sd1043/*1043:xpc10*/;
                       Tsf0SPILL10_256 <= 32'sd0;
                       end 
                      
                  13'sd1046/*1046:xpc10*/:  begin 
                       xpc10 <= 13'sd1047/*1047:xpc10*/;
                       Tsa1_SPILL_256 <= Tdsi1_5_V_0;
                       end 
                      
                  13'sd1050/*1050:xpc10*/: if (!(!Tsad1_3_V_1))  xpc10 <= 13'sd1294/*1294:xpc10*/;
                       else  xpc10 <= 13'sd1051/*1051:xpc10*/;

                  13'sd1054/*1054:xpc10*/:  begin 
                       xpc10 <= 13'sd1055/*1055:xpc10*/;
                       Tsad1_3_V_6 <= -32'sd1+Tsad1_3_V_6;
                       end 
                      
                  13'sd1058/*1058:xpc10*/: if (!(!rtl_signed_bitextract0(Tsad1_3_V_6)))  xpc10 <= 13'sd1253/*1253:xpc10*/;
                       else  xpc10 <= 13'sd1059/*1059:xpc10*/;

                  13'sd1062/*1062:xpc10*/:  begin 
                       xpc10 <= 13'sd1063/*1063:xpc10*/;
                       Tssh8_5_V_0 <= Tsad1_3_V_4;
                       end 
                      
                  13'sd1066/*1066:xpc10*/:  begin 
                       xpc10 <= 13'sd1067/*1067:xpc10*/;
                       Tsad1_3_V_4 <= Tssh8_5_V_0;
                       end 
                      
                  13'sd1067/*1067:xpc10*/:  begin 
                       xpc10 <= 13'sd1068/*1068:xpc10*/;
                       Tsad1_3_V_2 <= rtl_signed_bitextract0(Tsad1_3_V_0);
                       end 
                      
                  13'sd1071/*1071:xpc10*/:  begin 
                       xpc10 <= 13'sd1072/*1072:xpc10*/;
                       Tsad1_3_V_3 <= 64'sh_2000_0000_0000_0000|Tsad1_3_V_3;
                       end 
                      
                  13'sd1072/*1072:xpc10*/:  begin 
                       xpc10 <= 13'sd1073/*1073:xpc10*/;
                       Tsad1_3_V_5 <= (Tsad1_3_V_3+Tsad1_3_V_4<<32'sd1);
                       end 
                      
                  13'sd1073/*1073:xpc10*/:  begin 
                       xpc10 <= 13'sd1074/*1074:xpc10*/;
                       Tsad1_3_V_2 <= rtl_signed_bitextract0(-16'sd1+Tsad1_3_V_2);
                       end 
                      
                  13'sd1074/*1074:xpc10*/: if ((Tsad1_3_V_5<64'sh0))  xpc10 <= 13'sd1075/*1075:xpc10*/;
                       else  xpc10 <= 13'sd1081/*1081:xpc10*/;

                  13'sd1078/*1078:xpc10*/:  begin 
                       xpc10 <= 13'sd1079/*1079:xpc10*/;
                       Tsad1_3_V_5 <= Tsad1_3_V_3+Tsad1_3_V_4;
                       end 
                      
                  13'sd1079/*1079:xpc10*/:  begin 
                       xpc10 <= 13'sd1080/*1080:xpc10*/;
                       Tsad1_3_V_2 <= rtl_signed_bitextract0(16'sd1+Tsad1_3_V_2);
                       end 
                      
                  13'sd1083/*1083:xpc10*/:  begin 
                       xpc10 <= 13'sd1084/*1084:xpc10*/;
                       Tsro28_4_V_0 <= rtl_signed_bitextract0(Tsad1_3_V_2);
                       end 
                      
                  13'sd1084/*1084:xpc10*/:  begin 
                       xpc10 <= 13'sd1085/*1085:xpc10*/;
                       Tsro28_4_V_1 <= Tsad1_3_V_5;
                       end 
                      
                  13'sd1087/*1087:xpc10*/:  begin 
                       xpc10 <= 13'sd1088/*1088:xpc10*/;
                       Tsro28_4_V_5 <= 16'sh200;
                       end 
                      
                  13'sd1091/*1091:xpc10*/:  begin 
                       xpc10 <= 13'sd1092/*1092:xpc10*/;
                       Tsro28_4_V_6 <= rtl_signed_bitextract2(64'sh3ff&Tsro28_4_V_1);
                       end 
                      
                  13'sd1092/*1092:xpc10*/: if ((Tsro28_4_V_0<32'sd2045))  xpc10 <= 13'sd1171/*1171:xpc10*/;
                       else  xpc10 <= 13'sd1093/*1093:xpc10*/;

                  13'sd1096/*1096:xpc10*/: if ((32'sd2045<Tsro28_4_V_0))  xpc10 <= 13'sd1106/*1106:xpc10*/;
                       else  xpc10 <= 13'sd1097/*1097:xpc10*/;
              endcase
              if ((64'sh_3ee4_f8b5_88e3_68f1==(64'sh_7fff_ffff_ffff_ffff&Tdsi1_5_V_1)))  begin if ((13'sd998/*998:xpc10*/==xpc10))  xpc10
                       <= 13'sd1008/*1008:xpc10*/;

                       end 
                   else if ((13'sd998/*998:xpc10*/==xpc10))  xpc10 <= 13'sd999/*999:xpc10*/;
                      
              case (xpc10)
                  13'sd938/*938:xpc10*/:  xpc10 <= 13'sd939/*939:xpc10*/;

                  13'sd943/*943:xpc10*/:  xpc10 <= 13'sd944/*944:xpc10*/;

                  13'sd945/*945:xpc10*/:  begin 
                       xpc10 <= 13'sd946/*946:xpc10*/;
                       done <= 1'h1;
                       end 
                      
                  13'sd951/*951:xpc10*/:  xpc10 <= 13'sd952/*952:xpc10*/;

                  13'sd956/*956:xpc10*/:  begin 
                       xpc10 <= 13'sd957/*957:xpc10*/;
                       Tdb0_SPILL_258 <= 32'sd0;
                       end 
                      
                  13'sd957/*957:xpc10*/:  begin 
                       xpc10 <= 13'sd958/*958:xpc10*/;
                       Tdb0_SPILL_257 <= Tdb0_SPILL_259;
                       end 
                      
                  13'sd964/*964:xpc10*/:  begin 
                       xpc10 <= 13'sd965/*965:xpc10*/;
                       Tse5_SPILL_256 <= 32'sd0;
                       end 
                      
                  13'sd968/*968:xpc10*/:  begin 
                       xpc10 <= 13'sd969/*969:xpc10*/;
                       Tsfl0_3_V_0 <= rtl_unsigned_bitextract4(Tse5_SPILL_256);
                       end 
                      
                  13'sd969/*969:xpc10*/: if ((64'sh0<((64'sh_7fff_ffff_ffff_ffff&Tdsi1_5_V_1)>>32'sd63)))  xpc10 <= 13'sd970/*970:xpc10*/;
                       else  xpc10 <= 13'sd1012/*1012:xpc10*/;

                  13'sd973/*973:xpc10*/:  begin 
                       xpc10 <= 13'sd974/*974:xpc10*/;
                       Tse5SPILL10_256 <= 32'sd1;
                       end 
                      
                  13'sd977/*977:xpc10*/:  begin 
                       xpc10 <= 13'sd978/*978:xpc10*/;
                       Tsfl0_3_V_1 <= rtl_unsigned_bitextract4(Tse5SPILL10_256);
                       end 
                      
                  13'sd978/*978:xpc10*/:  begin 
                      if ((Tsfl0_3_V_0? !Tsfl0_3_V_1: Tsfl0_3_V_1))  begin if ((Tsfl0_3_V_0? !Tsfl0_3_V_1: Tsfl0_3_V_1))  xpc10 <= 13'sd979
                              /*979:xpc10*/;

                               end 
                          if ((Tsfl0_3_V_0? Tsfl0_3_V_1: !Tsfl0_3_V_1))  begin if ((Tsfl0_3_V_0? Tsfl0_3_V_1: !Tsfl0_3_V_1))  xpc10 <= 13'sd996
                              /*996:xpc10*/;

                               end 
                           end 
                      
                  13'sd982/*982:xpc10*/: if (Tsfl0_3_V_0)  xpc10 <= 13'sd992/*992:xpc10*/;
                       else  xpc10 <= 13'sd983/*983:xpc10*/;

                  13'sd986/*986:xpc10*/:  begin 
                       xpc10 <= 13'sd987/*987:xpc10*/;
                       Tsf0SPILL14_257 <= rtl_sign_extend3((32'sd0/*0:USA170*/==((64'sh_3ee4_f8b5_88e3_68f1|64'sh_7fff_ffff_ffff_ffff
                      &Tdsi1_5_V_1)<<32'sd1)));

                       end 
                      
                  13'sd990/*990:xpc10*/:  begin 
                       xpc10 <= 13'sd991/*991:xpc10*/;
                       Tsf0SPILL14_256 <= Tsf0SPILL14_257;
                       end 
                      
                  13'sd994/*994:xpc10*/:  begin 
                       xpc10 <= 13'sd995/*995:xpc10*/;
                       Tsf0SPILL14_257 <= 32'sd1;
                       end 
                      endcase
              if ((Tdbm0_3_V_0==32'sd36/*36:Tdbm0.3_V_0*/))  begin if ((13'sd934/*934:xpc10*/==xpc10))  xpc10 <= 13'sd935/*935:xpc10*/;
                       end 
                   else if ((13'sd934/*934:xpc10*/==xpc10))  xpc10 <= 13'sd949/*949:xpc10*/;
                      
              case (xpc10)
                  13'sd918/*918:xpc10*/:  xpc10 <= 13'sd919/*919:xpc10*/;

                  13'sd923/*923:xpc10*/:  begin 
                       xpc10 <= 13'sd924/*924:xpc10*/;
                       Tdbm0_3_V_1 <= 32'sd1+Tdbm0_3_V_1;
                       end 
                      
                  13'sd927/*927:xpc10*/: if ((Tdbm0_3_V_1<32'sd2))  xpc10 <= 13'sd422/*422:xpc10*/;
                       else  xpc10 <= 13'sd928/*928:xpc10*/;

                  13'sd932/*932:xpc10*/:  xpc10 <= 13'sd933/*933:xpc10*/;
              endcase
              if ((32'sd0/*0:USA176*/==(Tdbm0_3_V_2^A_64_US_CC_SCALbx10_ARA0[Tdbm0_3_V_1])))  begin if ((13'sd914/*914:xpc10*/==xpc10
                  ))  xpc10 <= 13'sd921/*921:xpc10*/;
                       end 
                   else if ((13'sd914/*914:xpc10*/==xpc10))  xpc10 <= 13'sd915/*915:xpc10*/;
                      
              case (xpc10)
                  13'sd905/*905:xpc10*/:  begin 
                       xpc10 <= 13'sd906/*906:xpc10*/;
                       Tdb0_SPILL_258 <= 32'sd1;
                       end 
                      
                  13'sd906/*906:xpc10*/:  begin 
                       xpc10 <= 13'sd907/*907:xpc10*/;
                       Tdb0_SPILL_257 <= Tdb0_SPILL_256;
                       end 
                      
                  13'sd910/*910:xpc10*/:  begin 
                       xpc10 <= 13'sd911/*911:xpc10*/;
                       Tdbm0_3_V_0 <= Tdb0_SPILL_258+Tdb0_SPILL_257;
                       end 
                      
                  13'sd912/*912:xpc10*/:  xpc10 <= 13'sd913/*913:xpc10*/;
              endcase
              if ((Tdbm0_3_V_2==A_64_US_CC_SCALbx10_ARA0[Tdbm0_3_V_1]))  begin if ((13'sd901/*901:xpc10*/==xpc10))  xpc10 <= 13'sd902
                      /*902:xpc10*/;

                       end 
                   else if ((13'sd901/*901:xpc10*/==xpc10))  xpc10 <= 13'sd954/*954:xpc10*/;
                      
              case (xpc10)
                  13'sd887/*887:xpc10*/:  begin 
                       xpc10 <= 13'sd888/*888:xpc10*/;
                       Tsf0SPILL14_256 <= 32'sd0;
                       end 
                      
                  13'sd891/*891:xpc10*/: if (!(!Tsf0SPILL14_256))  xpc10 <= 13'sd518/*518:xpc10*/;
                       else  xpc10 <= 13'sd892/*892:xpc10*/;

                  13'sd895/*895:xpc10*/:  begin 
                       xpc10 <= 13'sd896/*896:xpc10*/;
                       Tdbm0_3_V_2 <= Tdsi1_5_V_0;
                       end 
                      
                  13'sd898/*898:xpc10*/:  begin 
                       xpc10 <= 13'sd899/*899:xpc10*/;
                       fastspilldup88 <= Tdbm0_3_V_0;
                       end 
                      
                  13'sd899/*899:xpc10*/:  begin 
                       xpc10 <= 13'sd900/*900:xpc10*/;
                       Tdb0_SPILL_259 <= fastspilldup88;
                       end 
                      
                  13'sd900/*900:xpc10*/:  begin 
                       xpc10 <= 13'sd901/*901:xpc10*/;
                       Tdb0_SPILL_256 <= fastspilldup88;
                       end 
                      endcase
              if ((32'sd0/*0:USA168*/==(52'sd4503599627370495&Tdsi1_5_V_1)))  begin if ((13'sd882/*882:xpc10*/==xpc10))  xpc10 <= 13'sd959
                      /*959:xpc10*/;

                       end 
                   else if ((13'sd882/*882:xpc10*/==xpc10))  xpc10 <= 13'sd883/*883:xpc10*/;
                      if ((32'sd2047/*2047:USA166*/==rtl_signed_bitextract2(64'sh7ff&((64'sh_7fff_ffff_ffff_ffff&Tdsi1_5_V_1)>>32'sd52
              ))))  begin if ((13'sd878/*878:xpc10*/==xpc10))  xpc10 <= 13'sd879/*879:xpc10*/;
                       end 
                   else if ((13'sd878/*878:xpc10*/==xpc10))  xpc10 <= 13'sd959/*959:xpc10*/;
                      
              case (xpc10)
                  13'sd840/*840:xpc10*/:  begin 
                       xpc10 <= 13'sd841/*841:xpc10*/;
                       Tsf0SPILL12_256 <= rtl_sign_extend3((32'sd0/*0:USA88*/==(32'sd0/*0:USA86*/==(64'sh7_ffff_ffff_ffff&Tspr3_2_V_1
                      ))));

                       end 
                      
                  13'sd844/*844:xpc10*/:  begin 
                       xpc10 <= 13'sd845/*845:xpc10*/;
                       Tspr3_2_V_4 <= rtl_unsigned_bitextract4(Tsf0SPILL12_256);
                       end 
                      
                  13'sd845/*845:xpc10*/:  begin 
                       xpc10 <= 13'sd846/*846:xpc10*/;
                       Tspr3_2_V_0 <= 64'sh8_0000_0000_0000|Tspr3_2_V_0;
                       end 
                      
                  13'sd846/*846:xpc10*/:  begin 
                       xpc10 <= 13'sd847/*847:xpc10*/;
                       Tspr3_2_V_1 <= 64'sh8_0000_0000_0000|Tspr3_2_V_1;
                       end 
                      
                  13'sd847/*847:xpc10*/:  begin 
                      if (Tspr3_2_V_2 || Tspr3_2_V_4)  begin if (Tspr3_2_V_2 || Tspr3_2_V_4)  xpc10 <= 13'sd848/*848:xpc10*/;
                               end 
                          if (!Tspr3_2_V_2 && !Tspr3_2_V_4)  xpc10 <= 13'sd853/*853:xpc10*/;
                           end 
                      
                  13'sd855/*855:xpc10*/: if (Tspr3_2_V_4)  xpc10 <= 13'sd856/*856:xpc10*/;
                       else  xpc10 <= 13'sd1016/*1016:xpc10*/;

                  13'sd859/*859:xpc10*/:  begin 
                       xpc10 <= 13'sd860/*860:xpc10*/;
                       Tsp3_SPILL_256 <= Tspr3_2_V_1;
                       end 
                      
                  13'sd863/*863:xpc10*/:  begin 
                       xpc10 <= 13'sd864/*864:xpc10*/;
                       Tsa1_SPILL_256 <= Tsp3_SPILL_256;
                       end 
                      
                  13'sd867/*867:xpc10*/:  begin 
                       xpc10 <= 13'sd868/*868:xpc10*/;
                       Tsf1SPILL14_256 <= Tsa1_SPILL_256;
                       end 
                      
                  13'sd871/*871:xpc10*/:  begin 
                       xpc10 <= 13'sd872/*872:xpc10*/;
                       Tdsi1_5_V_0 <= Tsf1SPILL14_256;
                       end 
                      
                  13'sd872/*872:xpc10*/:  xpc10 <= 13'sd873/*873:xpc10*/;

                  13'sd874/*874:xpc10*/:  begin 
                       xpc10 <= 13'sd875/*875:xpc10*/;
                       Tdsi1_5_V_2 <= 32'sd1+Tdsi1_5_V_2;
                       end 
                      endcase
              if ((32'sd4094/*4094:USA84*/==(64'shfff&(Tspr3_2_V_1>>32'sd51))))  begin if ((13'sd836/*836:xpc10*/==xpc10))  xpc10 <= 13'sd837
                      /*837:xpc10*/;

                       end 
                   else if ((13'sd836/*836:xpc10*/==xpc10))  xpc10 <= 13'sd1036/*1036:xpc10*/;
                      
              case (xpc10)
                  13'sd830/*830:xpc10*/:  begin 
                       xpc10 <= 13'sd831/*831:xpc10*/;
                       Tsf0SPILL10_256 <= rtl_sign_extend3((32'sd0/*0:USA82*/==(32'sd0/*0:USA80*/==(64'sh7_ffff_ffff_ffff&Tspr3_2_V_0
                      ))));

                       end 
                      
                  13'sd834/*834:xpc10*/:  begin 
                       xpc10 <= 13'sd835/*835:xpc10*/;
                       Tspr3_2_V_2 <= rtl_unsigned_bitextract4(Tsf0SPILL10_256);
                       end 
                      
                  13'sd835/*835:xpc10*/:  begin 
                       xpc10 <= 13'sd836/*836:xpc10*/;
                       Tspr3_2_V_3 <= (32'sd0<rtl_sign_extend5(54'sd9007199254740992)+(Tspr3_2_V_1<<32'sd1));
                       end 
                      endcase
              if ((32'sd4094/*4094:USA78*/==(64'shfff&(Tspr3_2_V_0>>32'sd51))))  begin if ((13'sd826/*826:xpc10*/==xpc10))  xpc10 <= 13'sd827
                      /*827:xpc10*/;

                       end 
                   else if ((13'sd826/*826:xpc10*/==xpc10))  xpc10 <= 13'sd1040/*1040:xpc10*/;
                      
              case (xpc10)
                  13'sd755/*755:xpc10*/:  begin 
                       xpc10 <= 13'sd756/*756:xpc10*/;
                       Tsf0SPILL12_256 <= rtl_sign_extend3((32'sd0/*0:USA48*/==(32'sd0/*0:USA46*/==(64'sh7_ffff_ffff_ffff&Tspr2_2_V_1
                      ))));

                       end 
                      
                  13'sd759/*759:xpc10*/:  begin 
                       xpc10 <= 13'sd760/*760:xpc10*/;
                       Tspr2_2_V_4 <= rtl_unsigned_bitextract4(Tsf0SPILL12_256);
                       end 
                      
                  13'sd760/*760:xpc10*/:  begin 
                       xpc10 <= 13'sd761/*761:xpc10*/;
                       Tspr2_2_V_0 <= 64'sh8_0000_0000_0000|Tspr2_2_V_0;
                       end 
                      
                  13'sd761/*761:xpc10*/:  begin 
                       xpc10 <= 13'sd762/*762:xpc10*/;
                       Tspr2_2_V_1 <= 64'sh8_0000_0000_0000|Tspr2_2_V_1;
                       end 
                      
                  13'sd762/*762:xpc10*/:  begin 
                      if (Tspr2_2_V_2 || Tspr2_2_V_4)  begin if (Tspr2_2_V_2 || Tspr2_2_V_4)  xpc10 <= 13'sd763/*763:xpc10*/;
                               end 
                          if (!Tspr2_2_V_2 && !Tspr2_2_V_4)  xpc10 <= 13'sd768/*768:xpc10*/;
                           end 
                      
                  13'sd770/*770:xpc10*/: if (Tspr2_2_V_4)  xpc10 <= 13'sd771/*771:xpc10*/;
                       else  xpc10 <= 13'sd2260/*2260:xpc10*/;

                  13'sd774/*774:xpc10*/:  begin 
                       xpc10 <= 13'sd775/*775:xpc10*/;
                       Tsp2_SPILL_256 <= Tspr2_2_V_1;
                       end 
                      
                  13'sd778/*778:xpc10*/:  begin 
                       xpc10 <= 13'sd779/*779:xpc10*/;
                       Tsf1SPILL12_256 <= Tsp2_SPILL_256;
                       end 
                      
                  13'sd782/*782:xpc10*/:  begin 
                       xpc10 <= 13'sd783/*783:xpc10*/;
                       Tdsi1_5_V_1 <= Tsf1SPILL12_256;
                       end 
                      
                  13'sd783/*783:xpc10*/: if ((64'sh0<(Tdsi1_5_V_0>>32'sd63)))  xpc10 <= 13'sd784/*784:xpc10*/;
                       else  xpc10 <= 13'sd2256/*2256:xpc10*/;

                  13'sd787/*787:xpc10*/:  begin 
                       xpc10 <= 13'sd788/*788:xpc10*/;
                       Tse0SPILL16_256 <= 32'sd1;
                       end 
                      
                  13'sd791/*791:xpc10*/:  begin 
                       xpc10 <= 13'sd792/*792:xpc10*/;
                       Tsfl1_39_V_0 <= rtl_unsigned_bitextract4(Tse0SPILL16_256);
                       end 
                      
                  13'sd796/*796:xpc10*/:  begin 
                       xpc10 <= 13'sd797/*797:xpc10*/;
                       Tse0SPILL18_256 <= 32'sd1;
                       end 
                      
                  13'sd800/*800:xpc10*/:  begin 
                       xpc10 <= 13'sd801/*801:xpc10*/;
                       Tsfl1_39_V_1 <= rtl_unsigned_bitextract4(Tse0SPILL18_256);
                       end 
                      
                  13'sd801/*801:xpc10*/:  begin 
                      if ((Tsfl1_39_V_0? Tsfl1_39_V_1: !Tsfl1_39_V_1))  begin if ((Tsfl1_39_V_0? Tsfl1_39_V_1: !Tsfl1_39_V_1))  xpc10
                               <= 13'sd802/*802:xpc10*/;

                               end 
                          if ((Tsfl1_39_V_0? !Tsfl1_39_V_1: Tsfl1_39_V_1))  begin if ((Tsfl1_39_V_0? !Tsfl1_39_V_1: Tsfl1_39_V_1))  xpc10
                               <= 13'sd1575/*1575:xpc10*/;

                               end 
                           end 
                      
                  13'sd805/*805:xpc10*/:  begin 
                       xpc10 <= 13'sd806/*806:xpc10*/;
                       Tsad1_3_V_3 <= 64'shf_ffff_ffff_ffff&Tdsi1_5_V_0;
                       end 
                      
                  13'sd806/*806:xpc10*/:  begin 
                       xpc10 <= 13'sd807/*807:xpc10*/;
                       Tsad1_3_V_0 <= rtl_signed_bitextract2(64'sh7ff&(Tdsi1_5_V_0>>32'sd52));
                       end 
                      
                  13'sd807/*807:xpc10*/:  begin 
                       xpc10 <= 13'sd808/*808:xpc10*/;
                       Tsad1_3_V_4 <= 64'shf_ffff_ffff_ffff&Tdsi1_5_V_1;
                       end 
                      
                  13'sd808/*808:xpc10*/:  begin 
                       xpc10 <= 13'sd809/*809:xpc10*/;
                       Tsad1_3_V_1 <= rtl_signed_bitextract2(64'sh7ff&(Tdsi1_5_V_1>>32'sd52));
                       end 
                      
                  13'sd809/*809:xpc10*/:  begin 
                       xpc10 <= 13'sd810/*810:xpc10*/;
                       Tsad1_3_V_6 <= rtl_sign_extend9(Tsad1_3_V_0)+(0-Tsad1_3_V_1);
                       end 
                      
                  13'sd810/*810:xpc10*/:  begin 
                       xpc10 <= 13'sd811/*811:xpc10*/;
                       Tsad1_3_V_3 <= (Tsad1_3_V_3<<32'sd9);
                       end 
                      
                  13'sd811/*811:xpc10*/:  begin 
                       xpc10 <= 13'sd812/*812:xpc10*/;
                       Tsad1_3_V_4 <= (Tsad1_3_V_4<<32'sd9);
                       end 
                      
                  13'sd812/*812:xpc10*/: if ((32'sd0<Tsad1_3_V_6))  xpc10 <= 13'sd813/*813:xpc10*/;
                       else  xpc10 <= 13'sd1298/*1298:xpc10*/;

                  13'sd824/*824:xpc10*/:  begin 
                       xpc10 <= 13'sd825/*825:xpc10*/;
                       Tspr3_2_V_0 <= Tdsi1_5_V_0;
                       end 
                      
                  13'sd825/*825:xpc10*/:  begin 
                       xpc10 <= 13'sd826/*826:xpc10*/;
                       Tspr3_2_V_1 <= Tdsi1_5_V_1;
                       end 
                      endcase
              if ((32'sd4094/*4094:USA44*/==(64'shfff&(Tspr2_2_V_1>>32'sd51))))  begin if ((13'sd751/*751:xpc10*/==xpc10))  xpc10 <= 13'sd752
                      /*752:xpc10*/;

                       end 
                   else if ((13'sd751/*751:xpc10*/==xpc10))  xpc10 <= 13'sd2280/*2280:xpc10*/;
                      
              case (xpc10)
                  13'sd745/*745:xpc10*/:  begin 
                       xpc10 <= 13'sd746/*746:xpc10*/;
                       Tsf0SPILL10_256 <= rtl_sign_extend3((32'sd0/*0:USA42*/==(32'sd0/*0:USA40*/==(64'sh7_ffff_ffff_ffff&Tspr2_2_V_0
                      ))));

                       end 
                      
                  13'sd749/*749:xpc10*/:  begin 
                       xpc10 <= 13'sd750/*750:xpc10*/;
                       Tspr2_2_V_2 <= rtl_unsigned_bitextract4(Tsf0SPILL10_256);
                       end 
                      
                  13'sd750/*750:xpc10*/:  begin 
                       xpc10 <= 13'sd751/*751:xpc10*/;
                       Tspr2_2_V_3 <= (32'sd0<rtl_sign_extend5(54'sd9007199254740992)+(Tspr2_2_V_1<<32'sd1));
                       end 
                      endcase
              if ((32'sd4094/*4094:USA38*/==(64'shfff&(Tspr2_2_V_0>>32'sd51))))  begin if ((13'sd741/*741:xpc10*/==xpc10))  xpc10 <= 13'sd742
                      /*742:xpc10*/;

                       end 
                   else if ((13'sd741/*741:xpc10*/==xpc10))  xpc10 <= 13'sd2284/*2284:xpc10*/;
                      
              case (xpc10)
                  13'sd739/*739:xpc10*/:  begin 
                       xpc10 <= 13'sd740/*740:xpc10*/;
                       Tspr2_2_V_0 <= Tsf1SPILL10_256;
                       end 
                      
                  13'sd740/*740:xpc10*/:  begin 
                       xpc10 <= 13'sd741/*741:xpc10*/;
                       Tspr2_2_V_1 <= Tsi1SPILL10_256;
                       end 
                      endcase
              if ((Tsfl1_35_V_3==32'sd2047/*2047:Tsfl1.35_V_3*/))  begin if ((13'sd731/*731:xpc10*/==xpc10))  xpc10 <= 13'sd732/*732:xpc10*/;
                       end 
                   else if ((13'sd731/*731:xpc10*/==xpc10))  xpc10 <= 13'sd2388/*2388:xpc10*/;
                      
              case (xpc10)
                  13'sd657/*657:xpc10*/:  begin 
                       xpc10 <= 13'sd658/*658:xpc10*/;
                       Tspr4_3_V_0 <= Tdsi1_5_V_1;
                       end 
                      
                  13'sd658/*658:xpc10*/:  begin 
                       xpc10 <= 13'sd659/*659:xpc10*/;
                       Tspr4_3_V_1 <= Tdsi1_5_V_3;
                       end 
                      
                  13'sd663/*663:xpc10*/:  begin 
                       xpc10 <= 13'sd664/*664:xpc10*/;
                       Tsf0SPILL10_256 <= rtl_sign_extend3((32'sd0/*0:USA14*/==(32'sd0/*0:USA12*/==(64'sh7_ffff_ffff_ffff&Tspr4_3_V_0
                      ))));

                       end 
                      
                  13'sd667/*667:xpc10*/:  begin 
                       xpc10 <= 13'sd668/*668:xpc10*/;
                       Tspr4_3_V_2 <= rtl_unsigned_bitextract4(Tsf0SPILL10_256);
                       end 
                      
                  13'sd668/*668:xpc10*/:  begin 
                       xpc10 <= 13'sd669/*669:xpc10*/;
                       Tspr4_3_V_3 <= (32'sd0<rtl_sign_extend5(54'sd9007199254740992)+(Tspr4_3_V_1<<32'sd1));
                       end 
                      
                  13'sd673/*673:xpc10*/:  begin 
                       xpc10 <= 13'sd674/*674:xpc10*/;
                       Tsf0SPILL12_256 <= rtl_sign_extend3((32'sd0/*0:USA20*/==(32'sd0/*0:USA18*/==(64'sh7_ffff_ffff_ffff&Tspr4_3_V_1
                      ))));

                       end 
                      
                  13'sd677/*677:xpc10*/:  begin 
                       xpc10 <= 13'sd678/*678:xpc10*/;
                       Tspr4_3_V_4 <= rtl_unsigned_bitextract4(Tsf0SPILL12_256);
                       end 
                      
                  13'sd678/*678:xpc10*/:  begin 
                       xpc10 <= 13'sd679/*679:xpc10*/;
                       Tspr4_3_V_0 <= 64'sh8_0000_0000_0000|Tspr4_3_V_0;
                       end 
                      
                  13'sd679/*679:xpc10*/:  begin 
                       xpc10 <= 13'sd680/*680:xpc10*/;
                       Tspr4_3_V_1 <= 64'sh8_0000_0000_0000|Tspr4_3_V_1;
                       end 
                      
                  13'sd692/*692:xpc10*/:  begin 
                       xpc10 <= 13'sd693/*693:xpc10*/;
                       Tsp4_SPILL_256 <= Tspr4_3_V_1;
                       end 
                      
                  13'sd696/*696:xpc10*/:  begin 
                       xpc10 <= 13'sd697/*697:xpc10*/;
                       Tsf1SPILL10_256 <= Tsp4_SPILL_256;
                       end 
                      
                  13'sd704/*704:xpc10*/:  begin 
                       xpc10 <= 13'sd705/*705:xpc10*/;
                       Tsi1SPILL10_256 <= 64'h0;
                       end 
                      
                  13'sd708/*708:xpc10*/:  begin 
                       xpc10 <= 13'sd709/*709:xpc10*/;
                       Tsfl1_35_V_6 <= 64'shf_ffff_ffff_ffff&Tsf1SPILL10_256;
                       end 
                      
                  13'sd709/*709:xpc10*/:  begin 
                       xpc10 <= 13'sd710/*710:xpc10*/;
                       Tsfl1_35_V_3 <= rtl_signed_bitextract2(64'sh7ff&(Tsf1SPILL10_256>>32'sd52));
                       end 
                      
                  13'sd710/*710:xpc10*/: if ((64'sh0<(Tsf1SPILL10_256>>32'sd63)))  xpc10 <= 13'sd711/*711:xpc10*/;
                       else  xpc10 <= 13'sd3113/*3113:xpc10*/;

                  13'sd714/*714:xpc10*/:  begin 
                       xpc10 <= 13'sd715/*715:xpc10*/;
                       Tse0SPILL12_256 <= 32'sd1;
                       end 
                      
                  13'sd718/*718:xpc10*/:  begin 
                       xpc10 <= 13'sd719/*719:xpc10*/;
                       Tsfl1_35_V_0 <= rtl_unsigned_bitextract4(Tse0SPILL12_256);
                       end 
                      
                  13'sd719/*719:xpc10*/:  begin 
                       xpc10 <= 13'sd720/*720:xpc10*/;
                       Tsfl1_35_V_7 <= 64'shf_ffff_ffff_ffff&Tsi1SPILL10_256;
                       end 
                      
                  13'sd720/*720:xpc10*/:  begin 
                       xpc10 <= 13'sd721/*721:xpc10*/;
                       Tsfl1_35_V_4 <= rtl_signed_bitextract2(64'sh7ff&(Tsi1SPILL10_256>>32'sd52));
                       end 
                      
                  13'sd721/*721:xpc10*/: if ((64'sh0<(Tsi1SPILL10_256>>32'sd63)))  xpc10 <= 13'sd722/*722:xpc10*/;
                       else  xpc10 <= 13'sd3109/*3109:xpc10*/;

                  13'sd725/*725:xpc10*/:  begin 
                       xpc10 <= 13'sd726/*726:xpc10*/;
                       Tse0SPILL14_256 <= 32'sd1;
                       end 
                      
                  13'sd729/*729:xpc10*/:  begin 
                       xpc10 <= 13'sd730/*730:xpc10*/;
                       Tsfl1_35_V_1 <= rtl_unsigned_bitextract4(Tse0SPILL14_256);
                       end 
                      
                  13'sd730/*730:xpc10*/:  begin 
                       xpc10 <= 13'sd731/*731:xpc10*/;
                       Tsfl1_35_V_2 <= rtl_unsigned_bitextract12(Tsfl1_35_V_0^Tsfl1_35_V_1);
                       end 
                      endcase
              if ((Tsfl1_24_V_3==32'sd2047/*2047:Tsfl1.24_V_3*/))  begin if ((13'sd641/*641:xpc10*/==xpc10))  xpc10 <= 13'sd642/*642:xpc10*/;
                       end 
                   else if ((13'sd641/*641:xpc10*/==xpc10))  xpc10 <= 13'sd3227/*3227:xpc10*/;
                      
              case (xpc10)
                  13'sd563/*563:xpc10*/:  begin 
                       xpc10 <= 13'sd564/*564:xpc10*/;
                       Tspr4_3_V_0 <= Tdsi1_5_V_1;
                       end 
                      
                  13'sd564/*564:xpc10*/:  begin 
                       xpc10 <= 13'sd565/*565:xpc10*/;
                       Tspr4_3_V_1 <= Tdsi1_5_V_3;
                       end 
                      
                  13'sd569/*569:xpc10*/:  begin 
                       xpc10 <= 13'sd570/*570:xpc10*/;
                       Tsf0SPILL10_256 <= rtl_sign_extend3((32'sd0/*0:USA14*/==(32'sd0/*0:USA12*/==(64'sh7_ffff_ffff_ffff&Tspr4_3_V_0
                      ))));

                       end 
                      
                  13'sd573/*573:xpc10*/:  begin 
                       xpc10 <= 13'sd574/*574:xpc10*/;
                       Tspr4_3_V_2 <= rtl_unsigned_bitextract4(Tsf0SPILL10_256);
                       end 
                      
                  13'sd574/*574:xpc10*/:  begin 
                       xpc10 <= 13'sd575/*575:xpc10*/;
                       Tspr4_3_V_3 <= (32'sd0<rtl_sign_extend5(54'sd9007199254740992)+(Tspr4_3_V_1<<32'sd1));
                       end 
                      
                  13'sd579/*579:xpc10*/:  begin 
                       xpc10 <= 13'sd580/*580:xpc10*/;
                       Tsf0SPILL12_256 <= rtl_sign_extend3((32'sd0/*0:USA20*/==(32'sd0/*0:USA18*/==(64'sh7_ffff_ffff_ffff&Tspr4_3_V_1
                      ))));

                       end 
                      
                  13'sd583/*583:xpc10*/:  begin 
                       xpc10 <= 13'sd584/*584:xpc10*/;
                       Tspr4_3_V_4 <= rtl_unsigned_bitextract4(Tsf0SPILL12_256);
                       end 
                      
                  13'sd584/*584:xpc10*/:  begin 
                       xpc10 <= 13'sd585/*585:xpc10*/;
                       Tspr4_3_V_0 <= 64'sh8_0000_0000_0000|Tspr4_3_V_0;
                       end 
                      
                  13'sd585/*585:xpc10*/:  begin 
                       xpc10 <= 13'sd586/*586:xpc10*/;
                       Tspr4_3_V_1 <= 64'sh8_0000_0000_0000|Tspr4_3_V_1;
                       end 
                      
                  13'sd598/*598:xpc10*/:  begin 
                       xpc10 <= 13'sd599/*599:xpc10*/;
                       Tsp4_SPILL_256 <= Tspr4_3_V_1;
                       end 
                      
                  13'sd602/*602:xpc10*/:  begin 
                       xpc10 <= 13'sd603/*603:xpc10*/;
                       Tsf1_SPILL_256 <= Tsp4_SPILL_256;
                       end 
                      
                  13'sd610/*610:xpc10*/:  begin 
                       xpc10 <= 13'sd611/*611:xpc10*/;
                       Tsi1_SPILL_256 <= 64'h0;
                       end 
                      
                  13'sd614/*614:xpc10*/:  xpc10 <= 13'sd615/*615:xpc10*/;

                  13'sd616/*616:xpc10*/:  begin 
                       xpc10 <= 13'sd617/*617:xpc10*/;
                       Tsfl1_24_V_8 <= 64'h0;
                       end 
                      
                  13'sd617/*617:xpc10*/:  begin 
                       xpc10 <= 13'sd618/*618:xpc10*/;
                       Tsfl1_24_V_9 <= 64'h0;
                       end 
                      
                  13'sd618/*618:xpc10*/:  begin 
                       xpc10 <= 13'sd619/*619:xpc10*/;
                       Tsfl1_24_V_6 <= 64'shf_ffff_ffff_ffff&Tdsi1_5_V_1;
                       end 
                      
                  13'sd619/*619:xpc10*/:  begin 
                       xpc10 <= 13'sd620/*620:xpc10*/;
                       Tsfl1_24_V_3 <= rtl_signed_bitextract2(64'sh7ff&(Tdsi1_5_V_1>>32'sd52));
                       end 
                      
                  13'sd624/*624:xpc10*/:  begin 
                       xpc10 <= 13'sd625/*625:xpc10*/;
                       Tse0_SPILL_256 <= 32'sd1;
                       end 
                      
                  13'sd628/*628:xpc10*/:  begin 
                       xpc10 <= 13'sd629/*629:xpc10*/;
                       Tsfl1_24_V_0 <= rtl_unsigned_bitextract4(Tse0_SPILL_256);
                       end 
                      
                  13'sd629/*629:xpc10*/:  begin 
                       xpc10 <= 13'sd630/*630:xpc10*/;
                       Tsfl1_24_V_7 <= 64'shf_ffff_ffff_ffff&Tdsi1_5_V_3;
                       end 
                      
                  13'sd630/*630:xpc10*/:  begin 
                       xpc10 <= 13'sd631/*631:xpc10*/;
                       Tsfl1_24_V_4 <= rtl_signed_bitextract2(64'sh7ff&(Tdsi1_5_V_3>>32'sd52));
                       end 
                      
                  13'sd635/*635:xpc10*/:  begin 
                       xpc10 <= 13'sd636/*636:xpc10*/;
                       Tse0SPILL10_256 <= 32'sd1;
                       end 
                      
                  13'sd639/*639:xpc10*/:  begin 
                       xpc10 <= 13'sd640/*640:xpc10*/;
                       Tsfl1_24_V_1 <= rtl_unsigned_bitextract4(Tse0SPILL10_256);
                       end 
                      
                  13'sd640/*640:xpc10*/:  begin 
                       xpc10 <= 13'sd641/*641:xpc10*/;
                       Tsfl1_24_V_2 <= rtl_unsigned_bitextract12(Tsfl1_24_V_0^Tsfl1_24_V_1);
                       end 
                      endcase
              if ((Tsfl1_8_V_3==32'sd2047/*2047:Tsfl1.8_V_3*/))  begin if ((13'sd547/*547:xpc10*/==xpc10))  xpc10 <= 13'sd548/*548:xpc10*/;
                       end 
                   else if ((13'sd547/*547:xpc10*/==xpc10))  xpc10 <= 13'sd3849/*3849:xpc10*/;
                      
              case (xpc10)
                  13'sd470/*470:xpc10*/:  begin 
                       xpc10 <= 13'sd471/*471:xpc10*/;
                       Tspr4_3_V_0 <= $unsigned(A_64_US_CC_SCALbx12_ARB0[Tdbm0_3_V_1]);
                       end 
                      
                  13'sd471/*471:xpc10*/:  begin 
                       xpc10 <= 13'sd472/*472:xpc10*/;
                       Tspr4_3_V_1 <= $unsigned(A_64_US_CC_SCALbx12_ARB0[Tdbm0_3_V_1]);
                       end 
                      
                  13'sd476/*476:xpc10*/:  begin 
                       xpc10 <= 13'sd477/*477:xpc10*/;
                       Tsf0SPILL10_256 <= rtl_sign_extend3((32'sd0/*0:USA14*/==(32'sd0/*0:USA12*/==(64'sh7_ffff_ffff_ffff&Tspr4_3_V_0
                      ))));

                       end 
                      
                  13'sd480/*480:xpc10*/:  begin 
                       xpc10 <= 13'sd481/*481:xpc10*/;
                       Tspr4_3_V_2 <= rtl_unsigned_bitextract4(Tsf0SPILL10_256);
                       end 
                      
                  13'sd481/*481:xpc10*/:  begin 
                       xpc10 <= 13'sd482/*482:xpc10*/;
                       Tspr4_3_V_3 <= (32'sd0<rtl_sign_extend5(54'sd9007199254740992)+(Tspr4_3_V_1<<32'sd1));
                       end 
                      
                  13'sd486/*486:xpc10*/:  begin 
                       xpc10 <= 13'sd487/*487:xpc10*/;
                       Tsf0SPILL12_256 <= rtl_sign_extend3((32'sd0/*0:USA20*/==(32'sd0/*0:USA18*/==(64'sh7_ffff_ffff_ffff&Tspr4_3_V_1
                      ))));

                       end 
                      
                  13'sd490/*490:xpc10*/:  begin 
                       xpc10 <= 13'sd491/*491:xpc10*/;
                       Tspr4_3_V_4 <= rtl_unsigned_bitextract4(Tsf0SPILL12_256);
                       end 
                      
                  13'sd491/*491:xpc10*/:  begin 
                       xpc10 <= 13'sd492/*492:xpc10*/;
                       Tspr4_3_V_0 <= 64'sh8_0000_0000_0000|Tspr4_3_V_0;
                       end 
                      
                  13'sd492/*492:xpc10*/:  begin 
                       xpc10 <= 13'sd493/*493:xpc10*/;
                       Tspr4_3_V_1 <= 64'sh8_0000_0000_0000|Tspr4_3_V_1;
                       end 
                      
                  13'sd505/*505:xpc10*/:  begin 
                       xpc10 <= 13'sd506/*506:xpc10*/;
                       Tsp4_SPILL_256 <= Tspr4_3_V_1;
                       end 
                      
                  13'sd509/*509:xpc10*/:  begin 
                       xpc10 <= 13'sd510/*510:xpc10*/;
                       Tsf0_SPILL_256 <= Tsp4_SPILL_256;
                       end 
                      
                  13'sd513/*513:xpc10*/:  begin 
                       xpc10 <= 13'sd514/*514:xpc10*/;
                       Tsfl0_10_V_0 <= -64'sh_8000_0000_0000_0000&~Tsf0_SPILL_256|64'sh_7fff_ffff_ffff_ffff&Tsf0_SPILL_256;
                       end 
                      
                  13'sd514/*514:xpc10*/:  begin 
                       xpc10 <= 13'sd515/*515:xpc10*/;
                       Tdsi1_5_V_3 <= Tsfl0_10_V_0;
                       end 
                      
                  13'sd515/*515:xpc10*/:  xpc10 <= 13'sd516/*516:xpc10*/;

                  13'sd520/*520:xpc10*/:  xpc10 <= 13'sd521/*521:xpc10*/;

                  13'sd522/*522:xpc10*/:  begin 
                       xpc10 <= 13'sd523/*523:xpc10*/;
                       Tsfl1_8_V_8 <= 64'h0;
                       end 
                      
                  13'sd523/*523:xpc10*/:  begin 
                       xpc10 <= 13'sd524/*524:xpc10*/;
                       Tsfl1_8_V_9 <= 64'h0;
                       end 
                      
                  13'sd524/*524:xpc10*/:  begin 
                       xpc10 <= 13'sd525/*525:xpc10*/;
                       Tsfl1_8_V_6 <= 64'shf_ffff_ffff_ffff&Tdsi1_5_V_1;
                       end 
                      
                  13'sd525/*525:xpc10*/:  begin 
                       xpc10 <= 13'sd526/*526:xpc10*/;
                       Tsfl1_8_V_3 <= rtl_signed_bitextract2(64'sh7ff&(Tdsi1_5_V_1>>32'sd52));
                       end 
                      
                  13'sd530/*530:xpc10*/:  begin 
                       xpc10 <= 13'sd531/*531:xpc10*/;
                       Tse0_SPILL_256 <= 32'sd1;
                       end 
                      
                  13'sd534/*534:xpc10*/:  begin 
                       xpc10 <= 13'sd535/*535:xpc10*/;
                       Tsfl1_8_V_0 <= rtl_unsigned_bitextract4(Tse0_SPILL_256);
                       end 
                      
                  13'sd535/*535:xpc10*/:  begin 
                       xpc10 <= 13'sd536/*536:xpc10*/;
                       Tsfl1_8_V_7 <= 64'shf_ffff_ffff_ffff&Tdsi1_5_V_3;
                       end 
                      
                  13'sd536/*536:xpc10*/:  begin 
                       xpc10 <= 13'sd537/*537:xpc10*/;
                       Tsfl1_8_V_4 <= rtl_signed_bitextract2(64'sh7ff&(Tdsi1_5_V_3>>32'sd52));
                       end 
                      
                  13'sd541/*541:xpc10*/:  begin 
                       xpc10 <= 13'sd542/*542:xpc10*/;
                       Tse0SPILL10_256 <= 32'sd1;
                       end 
                      
                  13'sd545/*545:xpc10*/:  begin 
                       xpc10 <= 13'sd546/*546:xpc10*/;
                       Tsfl1_8_V_1 <= rtl_unsigned_bitextract4(Tse0SPILL10_256);
                       end 
                      
                  13'sd546/*546:xpc10*/:  begin 
                       xpc10 <= 13'sd547/*547:xpc10*/;
                       Tsfl1_8_V_2 <= rtl_unsigned_bitextract12(Tsfl1_8_V_0^Tsfl1_8_V_1);
                       end 
                      endcase
              if ((Tsfl0_9_V_3==32'sd2047/*2047:Tsfl0.9_V_3*/))  begin if ((13'sd454/*454:xpc10*/==xpc10))  xpc10 <= 13'sd455/*455:xpc10*/;
                       end 
                   else if ((13'sd454/*454:xpc10*/==xpc10))  xpc10 <= 13'sd4418/*4418:xpc10*/;
                      
              case (xpc10)
                  13'sd46/*46:xpc10*/:  begin 
                       xpc10 <= 13'sd47/*47:xpc10*/;
                       A_64_US_CC_SCALbx12_ARB0[64'd0] <= 64'd0;
                       end 
                      
                  13'sd47/*47:xpc10*/:  begin 
                       xpc10 <= 13'sd48/*48:xpc10*/;
                       A_64_US_CC_SCALbx12_ARB0[64'd1] <= 64'sh_3fc6_5717_fced_55c1;
                       end 
                      
                  13'sd48/*48:xpc10*/:  begin 
                       xpc10 <= 13'sd49/*49:xpc10*/;
                       A_64_US_CC_SCALbx12_ARB0[64'd2] <= 64'sh_3fd6_5717_fced_55c1;
                       end 
                      
                  13'sd49/*49:xpc10*/:  begin 
                       xpc10 <= 13'sd50/*50:xpc10*/;
                       A_64_US_CC_SCALbx12_ARB0[64'd3] <= 64'sh_3fe0_c151_fdb2_0051;
                       end 
                      
                  13'sd50/*50:xpc10*/:  begin 
                       xpc10 <= 13'sd51/*51:xpc10*/;
                       A_64_US_CC_SCALbx12_ARB0[64'd4] <= 64'sh_3fe6_5717_fced_55c1;
                       end 
                      
                  13'sd51/*51:xpc10*/:  begin 
                       xpc10 <= 13'sd52/*52:xpc10*/;
                       A_64_US_CC_SCALbx12_ARB0[64'd5] <= 64'sh_3feb_ecdd_fc28_ab31;
                       end 
                      
                  13'sd52/*52:xpc10*/:  begin 
                       xpc10 <= 13'sd53/*53:xpc10*/;
                       A_64_US_CC_SCALbx12_ARB0[64'd6] <= 64'sh_3ff0_c151_fdb2_0051;
                       end 
                      
                  13'sd53/*53:xpc10*/:  begin 
                       xpc10 <= 13'sd54/*54:xpc10*/;
                       A_64_US_CC_SCALbx12_ARB0[64'd7] <= 64'sh_3ff3_8c34_fd4f_ab09;
                       end 
                      
                  13'sd54/*54:xpc10*/:  begin 
                       xpc10 <= 13'sd55/*55:xpc10*/;
                       A_64_US_CC_SCALbx12_ARB0[64'd8] <= 64'sh_3ff6_5717_fced_55c1;
                       end 
                      
                  13'sd55/*55:xpc10*/:  begin 
                       xpc10 <= 13'sd56/*56:xpc10*/;
                       A_64_US_CC_SCALbx12_ARB0[64'd9] <= 64'sh_3ff9_21fa_fc8b_0079;
                       end 
                      
                  13'sd56/*56:xpc10*/:  begin 
                       xpc10 <= 13'sd57/*57:xpc10*/;
                       A_64_US_CC_SCALbx12_ARB0[64'd10] <= 64'sh_3ffb_ecdd_fc28_ab31;
                       end 
                      
                  13'sd57/*57:xpc10*/:  begin 
                       xpc10 <= 13'sd58/*58:xpc10*/;
                       A_64_US_CC_SCALbx12_ARB0[64'd11] <= 64'sh_3ffe_b7c0_fbc6_55e9;
                       end 
                      
                  13'sd58/*58:xpc10*/:  begin 
                       xpc10 <= 13'sd59/*59:xpc10*/;
                       A_64_US_CC_SCALbx12_ARB0[64'd12] <= 64'sh_4000_c151_fdb2_0051;
                       end 
                      
                  13'sd59/*59:xpc10*/:  begin 
                       xpc10 <= 13'sd60/*60:xpc10*/;
                       A_64_US_CC_SCALbx12_ARB0[64'd13] <= 64'sh_4002_26c3_7d80_d5ad;
                       end 
                      
                  13'sd60/*60:xpc10*/:  begin 
                       xpc10 <= 13'sd61/*61:xpc10*/;
                       A_64_US_CC_SCALbx12_ARB0[64'd14] <= 64'sh_4003_8c34_fd4f_ab09;
                       end 
                      
                  13'sd61/*61:xpc10*/:  begin 
                       xpc10 <= 13'sd62/*62:xpc10*/;
                       A_64_US_CC_SCALbx12_ARB0[64'd15] <= 64'sh_4004_f1a6_7d1e_8065;
                       end 
                      
                  13'sd62/*62:xpc10*/:  begin 
                       xpc10 <= 13'sd63/*63:xpc10*/;
                       A_64_US_CC_SCALbx12_ARB0[64'd16] <= 64'sh_4006_5717_fced_55c1;
                       end 
                      
                  13'sd63/*63:xpc10*/:  begin 
                       xpc10 <= 13'sd64/*64:xpc10*/;
                       A_64_US_CC_SCALbx12_ARB0[64'd17] <= 64'sh_4007_bc89_7cbc_2b1d;
                       end 
                      
                  13'sd64/*64:xpc10*/:  begin 
                       xpc10 <= 13'sd65/*65:xpc10*/;
                       A_64_US_CC_SCALbx12_ARB0[64'd18] <= 64'sh_4009_21fa_fc8b_0079;
                       end 
                      
                  13'sd65/*65:xpc10*/:  begin 
                       xpc10 <= 13'sd66/*66:xpc10*/;
                       A_64_US_CC_SCALbx12_ARB0[64'd19] <= 64'sh_400a_876c_7c59_d5d5;
                       end 
                      
                  13'sd66/*66:xpc10*/:  begin 
                       xpc10 <= 13'sd67/*67:xpc10*/;
                       A_64_US_CC_SCALbx12_ARB0[64'd20] <= 64'sh_400b_ecdd_fc28_ab31;
                       end 
                      
                  13'sd67/*67:xpc10*/:  begin 
                       xpc10 <= 13'sd68/*68:xpc10*/;
                       A_64_US_CC_SCALbx12_ARB0[64'd21] <= 64'sh_400d_524f_7bf7_808d;
                       end 
                      
                  13'sd68/*68:xpc10*/:  begin 
                       xpc10 <= 13'sd69/*69:xpc10*/;
                       A_64_US_CC_SCALbx12_ARB0[64'd22] <= 64'sh_400e_b7c0_fbc6_55e9;
                       end 
                      
                  13'sd69/*69:xpc10*/:  begin 
                       xpc10 <= 13'sd70/*70:xpc10*/;
                       A_64_US_CC_SCALbx12_ARB0[64'd23] <= 64'sh_4010_0e99_3dca_95a3;
                       end 
                      
                  13'sd70/*70:xpc10*/:  begin 
                       xpc10 <= 13'sd71/*71:xpc10*/;
                       A_64_US_CC_SCALbx12_ARB0[64'd24] <= 64'sh_4010_c151_fdb2_0051;
                       end 
                      
                  13'sd71/*71:xpc10*/:  begin 
                       xpc10 <= 13'sd72/*72:xpc10*/;
                       A_64_US_CC_SCALbx12_ARB0[64'd25] <= 64'sh_4011_740a_bd99_6aff;
                       end 
                      
                  13'sd72/*72:xpc10*/:  begin 
                       xpc10 <= 13'sd73/*73:xpc10*/;
                       A_64_US_CC_SCALbx12_ARB0[64'd26] <= 64'sh_4012_26c3_7d80_d5ad;
                       end 
                      
                  13'sd73/*73:xpc10*/:  begin 
                       xpc10 <= 13'sd74/*74:xpc10*/;
                       A_64_US_CC_SCALbx12_ARB0[64'd27] <= 64'sh_4012_d97c_3d68_405b;
                       end 
                      
                  13'sd74/*74:xpc10*/:  begin 
                       xpc10 <= 13'sd75/*75:xpc10*/;
                       A_64_US_CC_SCALbx12_ARB0[64'd28] <= 64'sh_4013_8c34_fd4f_ab09;
                       end 
                      
                  13'sd75/*75:xpc10*/:  begin 
                       xpc10 <= 13'sd76/*76:xpc10*/;
                       A_64_US_CC_SCALbx12_ARB0[64'd29] <= 64'sh_4014_3eed_bd37_15b7;
                       end 
                      
                  13'sd76/*76:xpc10*/:  begin 
                       xpc10 <= 13'sd77/*77:xpc10*/;
                       A_64_US_CC_SCALbx12_ARB0[64'd30] <= 64'sh_4014_f1a6_7d1e_8065;
                       end 
                      
                  13'sd77/*77:xpc10*/:  begin 
                       xpc10 <= 13'sd78/*78:xpc10*/;
                       A_64_US_CC_SCALbx12_ARB0[64'd31] <= 64'sh_4015_a45f_3d05_eb13;
                       end 
                      
                  13'sd78/*78:xpc10*/:  begin 
                       xpc10 <= 13'sd79/*79:xpc10*/;
                       A_64_US_CC_SCALbx12_ARB0[64'd32] <= 64'sh_4016_5717_fced_55c1;
                       end 
                      
                  13'sd79/*79:xpc10*/:  begin 
                       xpc10 <= 13'sd80/*80:xpc10*/;
                       A_64_US_CC_SCALbx12_ARB0[64'd33] <= 64'sh_4017_09d0_bcd4_c06f;
                       end 
                      
                  13'sd80/*80:xpc10*/:  begin 
                       xpc10 <= 13'sd81/*81:xpc10*/;
                       A_64_US_CC_SCALbx12_ARB0[64'd34] <= 64'sh_4017_bc89_7cbc_2b1d;
                       end 
                      
                  13'sd81/*81:xpc10*/:  begin 
                       xpc10 <= 13'sd82/*82:xpc10*/;
                       A_64_US_CC_SCALbx12_ARB0[64'd35] <= 64'sh_4018_6f42_3ca3_95cb;
                       end 
                      
                  13'sd85/*85:xpc10*/:  begin 
                       xpc10 <= 13'sd86/*86:xpc10*/;
                       A_64_US_CC_SCALbx10_ARA0[64'd0] <= 64'd0;
                       end 
                      
                  13'sd86/*86:xpc10*/:  begin 
                       xpc10 <= 13'sd87/*87:xpc10*/;
                       A_64_US_CC_SCALbx10_ARA0[64'd1] <= 64'sh_3fc6_3a1a_335a_adcd;
                       end 
                      
                  13'sd87/*87:xpc10*/:  begin 
                       xpc10 <= 13'sd88/*88:xpc10*/;
                       A_64_US_CC_SCALbx10_ARA0[64'd2] <= 64'sh_3fd5_e3a8_2b09_bf3e;
                       end 
                      
                  13'sd88/*88:xpc10*/:  begin 
                       xpc10 <= 13'sd89/*89:xpc10*/;
                       A_64_US_CC_SCALbx10_ARA0[64'd3] <= 64'sh_3fdf_ffff_91f9_aa91;
                       end 
                      
                  13'sd89/*89:xpc10*/:  begin 
                       xpc10 <= 13'sd90/*90:xpc10*/;
                       A_64_US_CC_SCALbx10_ARA0[64'd4] <= 64'sh_3fe4_91b7_16c2_42e3;
                       end 
                      
                  13'sd90/*90:xpc10*/:  begin 
                       xpc10 <= 13'sd91/*91:xpc10*/;
                       A_64_US_CC_SCALbx10_ARA0[64'd5] <= 64'sh_3fe8_836f_6726_14a6;
                       end 
                      
                  13'sd91/*91:xpc10*/:  begin 
                       xpc10 <= 13'sd92/*92:xpc10*/;
                       A_64_US_CC_SCALbx10_ARA0[64'd6] <= 64'sh_3feb_b67a_c40b_2bed;
                       end 
                      
                  13'sd92/*92:xpc10*/:  begin 
                       xpc10 <= 13'sd93/*93:xpc10*/;
                       A_64_US_CC_SCALbx10_ARA0[64'd7] <= 64'sh_3fee_11f6_127e_28ad;
                       end 
                      
                  13'sd93/*93:xpc10*/:  begin 
                       xpc10 <= 13'sd94/*94:xpc10*/;
                       A_64_US_CC_SCALbx10_ARA0[64'd8] <= 64'sh_3fef_838b_6adf_fac0;
                       end 
                      
                  13'sd94/*94:xpc10*/:  begin 
                       xpc10 <= 13'sd95/*95:xpc10*/;
                       A_64_US_CC_SCALbx10_ARA0[64'd9] <= 64'sh_3fef_ffff_e1cb_d7aa;
                       end 
                      
                  13'sd95/*95:xpc10*/:  begin 
                       xpc10 <= 13'sd96/*96:xpc10*/;
                       A_64_US_CC_SCALbx10_ARA0[64'd10] <= 64'sh_3fef_838b_b014_7989;
                       end 
                      
                  13'sd96/*96:xpc10*/:  begin 
                       xpc10 <= 13'sd97/*97:xpc10*/;
                       A_64_US_CC_SCALbx10_ARA0[64'd11] <= 64'sh_3fee_11f6_92d9_62b4;
                       end 
                      
                  13'sd97/*97:xpc10*/:  begin 
                       xpc10 <= 13'sd98/*98:xpc10*/;
                       A_64_US_CC_SCALbx10_ARA0[64'd12] <= 64'sh_3feb_b67b_77c0_142d;
                       end 
                      
                  13'sd98/*98:xpc10*/:  begin 
                       xpc10 <= 13'sd99/*99:xpc10*/;
                       A_64_US_CC_SCALbx10_ARA0[64'd13] <= 64'sh_3fe8_8370_9d4e_a869;
                       end 
                      
                  13'sd99/*99:xpc10*/:  begin 
                       xpc10 <= 13'sd100/*100:xpc10*/;
                       A_64_US_CC_SCALbx10_ARA0[64'd14] <= 64'sh_3fe4_91b8_1d72_d8e8;
                       end 
                      
                  13'sd100/*100:xpc10*/:  begin 
                       xpc10 <= 13'sd101/*101:xpc10*/;
                       A_64_US_CC_SCALbx10_ARA0[64'd15] <= 64'sh_3fe0_0000_ea5f_43c8;
                       end 
                      
                  13'sd101/*101:xpc10*/:  begin 
                       xpc10 <= 13'sd102/*102:xpc10*/;
                       A_64_US_CC_SCALbx10_ARA0[64'd16] <= 64'sh_3fd5_e3aa_4e05_90c5;
                       end 
                      
                  13'sd102/*102:xpc10*/:  begin 
                       xpc10 <= 13'sd103/*103:xpc10*/;
                       A_64_US_CC_SCALbx10_ARA0[64'd17] <= 64'sh_3fc6_3a1d_2189_552c;
                       end 
                      
                  13'sd103/*103:xpc10*/:  begin 
                       xpc10 <= 13'sd104/*104:xpc10*/;
                       A_64_US_CC_SCALbx10_ARA0[64'd18] <= 64'sh_3ea6_aedf_fc45_4b91;
                       end 
                      
                  13'sd104/*104:xpc10*/:  begin 
                       xpc10 <= 13'sd105/*105:xpc10*/;
                       A_64_US_CC_SCALbx10_ARA0[64'd19] <= -64'sh_4039_c5eb_bb22_4c84;
                       end 
                      
                  13'sd105/*105:xpc10*/:  begin 
                       xpc10 <= 13'sd106/*106:xpc10*/;
                       A_64_US_CC_SCALbx10_ARA0[64'd20] <= -64'sh_402a_1c5b_1970_70c2;
                       end 
                      
                  13'sd106/*106:xpc10*/:  begin 
                       xpc10 <= 13'sd107/*107:xpc10*/;
                       A_64_US_CC_SCALbx10_ARA0[64'd21] <= -64'sh_4020_0002_b6b3_0695;
                       end 
                      
                  13'sd107/*107:xpc10*/:  begin 
                       xpc10 <= 13'sd108/*108:xpc10*/;
                       A_64_US_CC_SCALbx10_ARA0[64'd22] <= -64'sh_401b_6e49_e346_5c2d;
                       end 
                      
                  13'sd108/*108:xpc10*/:  begin 
                       xpc10 <= 13'sd109/*109:xpc10*/;
                       A_64_US_CC_SCALbx10_ARA0[64'd23] <= -64'sh_4017_7c91_4d23_07eb;
                       end 
                      
                  13'sd109/*109:xpc10*/:  begin 
                       xpc10 <= 13'sd110/*110:xpc10*/;
                       A_64_US_CC_SCALbx10_ARA0[64'd24] <= -64'sh_4014_4985_8bf5_51ce;
                       end 
                      
                  13'sd110/*110:xpc10*/:  begin 
                       xpc10 <= 13'sd111/*111:xpc10*/;
                       A_64_US_CC_SCALbx10_ARA0[64'd25] <= -64'sh_4011_ee0a_6ed2_dea9;
                       end 
                      
                  13'sd111/*111:xpc10*/:  begin 
                       xpc10 <= 13'sd112/*112:xpc10*/;
                       A_64_US_CC_SCALbx10_ARA0[64'd26] <= -64'sh_4010_7c74_e539_b504;
                       end 
                      
                  13'sd112/*112:xpc10*/:  begin 
                       xpc10 <= 13'sd113/*113:xpc10*/;
                       A_64_US_CC_SCALbx10_ARA0[64'd27] <= -64'sh_4010_0000_3d1a_2371;
                       end 
                      
                  13'sd113/*113:xpc10*/:  begin 
                       xpc10 <= 13'sd114/*114:xpc10*/;
                       A_64_US_CC_SCALbx10_ARA0[64'd28] <= -64'sh_4010_7c74_a15d_1816;
                       end 
                      
                  13'sd114/*114:xpc10*/:  begin 
                       xpc10 <= 13'sd115/*115:xpc10*/;
                       A_64_US_CC_SCALbx10_ARA0[64'd29] <= -64'sh_4011_ee08_eed2_51d9;
                       end 
                      
                  13'sd115/*115:xpc10*/:  begin 
                       xpc10 <= 13'sd116/*116:xpc10*/;
                       A_64_US_CC_SCALbx10_ARA0[64'd30] <= -64'sh_4014_4983_d3ce_34b6;
                       end 
                      
                  13'sd116/*116:xpc10*/:  begin 
                       xpc10 <= 13'sd117/*117:xpc10*/;
                       A_64_US_CC_SCALbx10_ARA0[64'd31] <= -64'sh_4017_7c8e_9190_287f;
                       end 
                      
                  13'sd117/*117:xpc10*/:  begin 
                       xpc10 <= 13'sd118/*118:xpc10*/;
                       A_64_US_CC_SCALbx10_ARA0[64'd32] <= -64'sh_401b_6e46_32e4_a2aa;
                       end 
                      
                  13'sd118/*118:xpc10*/:  begin 
                       xpc10 <= 13'sd119/*119:xpc10*/;
                       A_64_US_CC_SCALbx10_ARA0[64'd33] <= -64'sh_401f_fffd_e2f3_5cf3;
                       end 
                      
                  13'sd119/*119:xpc10*/:  begin 
                       xpc10 <= 13'sd120/*120:xpc10*/;
                       A_64_US_CC_SCALbx10_ARA0[64'd34] <= -64'sh_402a_1c52_f596_3509;
                       end 
                      
                  13'sd120/*120:xpc10*/:  begin 
                       xpc10 <= 13'sd121/*121:xpc10*/;
                       A_64_US_CC_SCALbx10_ARA0[64'd35] <= -64'sh_4039_c5dc_3b77_9c23;
                       end 
                      
                  13'sd122/*122:xpc10*/:  begin 
                       xpc10 <= 13'sd123/*123:xpc10*/;
                       done <= 1'h0;
                       end 
                      
                  13'sd134/*134:xpc10*/:  begin 
                       xpc10 <= 13'sd135/*135:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[32'd0] <= 8'h8;
                       end 
                      
                  13'sd135/*135:xpc10*/:  begin 
                       xpc10 <= 13'sd136/*136:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh1] <= 8'h7;
                       end 
                      
                  13'sd136/*136:xpc10*/:  begin 
                       xpc10 <= 13'sd137/*137:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh2] <= 8'h6;
                       end 
                      
                  13'sd137/*137:xpc10*/:  begin 
                       xpc10 <= 13'sd138/*138:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh3] <= 8'h6;
                       end 
                      
                  13'sd138/*138:xpc10*/:  begin 
                       xpc10 <= 13'sd139/*139:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh4] <= 8'h5;
                       end 
                      
                  13'sd139/*139:xpc10*/:  begin 
                       xpc10 <= 13'sd140/*140:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh5] <= 8'h5;
                       end 
                      
                  13'sd140/*140:xpc10*/:  begin 
                       xpc10 <= 13'sd141/*141:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh6] <= 8'h5;
                       end 
                      
                  13'sd141/*141:xpc10*/:  begin 
                       xpc10 <= 13'sd142/*142:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh7] <= 8'h5;
                       end 
                      
                  13'sd142/*142:xpc10*/:  begin 
                       xpc10 <= 13'sd143/*143:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh8] <= 8'h4;
                       end 
                      
                  13'sd143/*143:xpc10*/:  begin 
                       xpc10 <= 13'sd144/*144:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh9] <= 8'h4;
                       end 
                      
                  13'sd144/*144:xpc10*/:  begin 
                       xpc10 <= 13'sd145/*145:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sha] <= 8'h4;
                       end 
                      
                  13'sd145/*145:xpc10*/:  begin 
                       xpc10 <= 13'sd146/*146:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shb] <= 8'h4;
                       end 
                      
                  13'sd146/*146:xpc10*/:  begin 
                       xpc10 <= 13'sd147/*147:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shc] <= 8'h4;
                       end 
                      
                  13'sd147/*147:xpc10*/:  begin 
                       xpc10 <= 13'sd148/*148:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shd] <= 8'h4;
                       end 
                      
                  13'sd148/*148:xpc10*/:  begin 
                       xpc10 <= 13'sd149/*149:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'she] <= 8'h4;
                       end 
                      
                  13'sd149/*149:xpc10*/:  begin 
                       xpc10 <= 13'sd150/*150:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shf] <= 8'h4;
                       end 
                      
                  13'sd150/*150:xpc10*/:  begin 
                       xpc10 <= 13'sd151/*151:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh10] <= 8'h3;
                       end 
                      
                  13'sd151/*151:xpc10*/:  begin 
                       xpc10 <= 13'sd152/*152:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh11] <= 8'h3;
                       end 
                      
                  13'sd152/*152:xpc10*/:  begin 
                       xpc10 <= 13'sd153/*153:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh12] <= 8'h3;
                       end 
                      
                  13'sd153/*153:xpc10*/:  begin 
                       xpc10 <= 13'sd154/*154:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh13] <= 8'h3;
                       end 
                      
                  13'sd154/*154:xpc10*/:  begin 
                       xpc10 <= 13'sd155/*155:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh14] <= 8'h3;
                       end 
                      
                  13'sd155/*155:xpc10*/:  begin 
                       xpc10 <= 13'sd156/*156:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh15] <= 8'h3;
                       end 
                      
                  13'sd156/*156:xpc10*/:  begin 
                       xpc10 <= 13'sd157/*157:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh16] <= 8'h3;
                       end 
                      
                  13'sd157/*157:xpc10*/:  begin 
                       xpc10 <= 13'sd158/*158:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh17] <= 8'h3;
                       end 
                      
                  13'sd158/*158:xpc10*/:  begin 
                       xpc10 <= 13'sd159/*159:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh18] <= 8'h3;
                       end 
                      
                  13'sd159/*159:xpc10*/:  begin 
                       xpc10 <= 13'sd160/*160:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh19] <= 8'h3;
                       end 
                      
                  13'sd160/*160:xpc10*/:  begin 
                       xpc10 <= 13'sd161/*161:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh1a] <= 8'h3;
                       end 
                      
                  13'sd161/*161:xpc10*/:  begin 
                       xpc10 <= 13'sd162/*162:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh1b] <= 8'h3;
                       end 
                      
                  13'sd162/*162:xpc10*/:  begin 
                       xpc10 <= 13'sd163/*163:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh1c] <= 8'h3;
                       end 
                      
                  13'sd163/*163:xpc10*/:  begin 
                       xpc10 <= 13'sd164/*164:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh1d] <= 8'h3;
                       end 
                      
                  13'sd164/*164:xpc10*/:  begin 
                       xpc10 <= 13'sd165/*165:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh1e] <= 8'h3;
                       end 
                      
                  13'sd165/*165:xpc10*/:  begin 
                       xpc10 <= 13'sd166/*166:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh1f] <= 8'h3;
                       end 
                      
                  13'sd166/*166:xpc10*/:  begin 
                       xpc10 <= 13'sd167/*167:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh20] <= 8'h2;
                       end 
                      
                  13'sd167/*167:xpc10*/:  begin 
                       xpc10 <= 13'sd168/*168:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh21] <= 8'h2;
                       end 
                      
                  13'sd168/*168:xpc10*/:  begin 
                       xpc10 <= 13'sd169/*169:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh22] <= 8'h2;
                       end 
                      
                  13'sd169/*169:xpc10*/:  begin 
                       xpc10 <= 13'sd170/*170:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh23] <= 8'h2;
                       end 
                      
                  13'sd170/*170:xpc10*/:  begin 
                       xpc10 <= 13'sd171/*171:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh24] <= 8'h2;
                       end 
                      
                  13'sd171/*171:xpc10*/:  begin 
                       xpc10 <= 13'sd172/*172:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh25] <= 8'h2;
                       end 
                      
                  13'sd172/*172:xpc10*/:  begin 
                       xpc10 <= 13'sd173/*173:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh26] <= 8'h2;
                       end 
                      
                  13'sd173/*173:xpc10*/:  begin 
                       xpc10 <= 13'sd174/*174:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh27] <= 8'h2;
                       end 
                      
                  13'sd174/*174:xpc10*/:  begin 
                       xpc10 <= 13'sd175/*175:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh28] <= 8'h2;
                       end 
                      
                  13'sd175/*175:xpc10*/:  begin 
                       xpc10 <= 13'sd176/*176:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh29] <= 8'h2;
                       end 
                      
                  13'sd176/*176:xpc10*/:  begin 
                       xpc10 <= 13'sd177/*177:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh2a] <= 8'h2;
                       end 
                      
                  13'sd177/*177:xpc10*/:  begin 
                       xpc10 <= 13'sd178/*178:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh2b] <= 8'h2;
                       end 
                      
                  13'sd178/*178:xpc10*/:  begin 
                       xpc10 <= 13'sd179/*179:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh2c] <= 8'h2;
                       end 
                      
                  13'sd179/*179:xpc10*/:  begin 
                       xpc10 <= 13'sd180/*180:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh2d] <= 8'h2;
                       end 
                      
                  13'sd180/*180:xpc10*/:  begin 
                       xpc10 <= 13'sd181/*181:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh2e] <= 8'h2;
                       end 
                      
                  13'sd181/*181:xpc10*/:  begin 
                       xpc10 <= 13'sd182/*182:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh2f] <= 8'h2;
                       end 
                      
                  13'sd182/*182:xpc10*/:  begin 
                       xpc10 <= 13'sd183/*183:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh30] <= 8'h2;
                       end 
                      
                  13'sd183/*183:xpc10*/:  begin 
                       xpc10 <= 13'sd184/*184:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh31] <= 8'h2;
                       end 
                      
                  13'sd184/*184:xpc10*/:  begin 
                       xpc10 <= 13'sd185/*185:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh32] <= 8'h2;
                       end 
                      
                  13'sd185/*185:xpc10*/:  begin 
                       xpc10 <= 13'sd186/*186:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh33] <= 8'h2;
                       end 
                      
                  13'sd186/*186:xpc10*/:  begin 
                       xpc10 <= 13'sd187/*187:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh34] <= 8'h2;
                       end 
                      
                  13'sd187/*187:xpc10*/:  begin 
                       xpc10 <= 13'sd188/*188:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh35] <= 8'h2;
                       end 
                      
                  13'sd188/*188:xpc10*/:  begin 
                       xpc10 <= 13'sd189/*189:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh36] <= 8'h2;
                       end 
                      
                  13'sd189/*189:xpc10*/:  begin 
                       xpc10 <= 13'sd190/*190:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh37] <= 8'h2;
                       end 
                      
                  13'sd190/*190:xpc10*/:  begin 
                       xpc10 <= 13'sd191/*191:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh38] <= 8'h2;
                       end 
                      
                  13'sd191/*191:xpc10*/:  begin 
                       xpc10 <= 13'sd192/*192:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh39] <= 8'h2;
                       end 
                      
                  13'sd192/*192:xpc10*/:  begin 
                       xpc10 <= 13'sd193/*193:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh3a] <= 8'h2;
                       end 
                      
                  13'sd193/*193:xpc10*/:  begin 
                       xpc10 <= 13'sd194/*194:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh3b] <= 8'h2;
                       end 
                      
                  13'sd194/*194:xpc10*/:  begin 
                       xpc10 <= 13'sd195/*195:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh3c] <= 8'h2;
                       end 
                      
                  13'sd195/*195:xpc10*/:  begin 
                       xpc10 <= 13'sd196/*196:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh3d] <= 8'h2;
                       end 
                      
                  13'sd196/*196:xpc10*/:  begin 
                       xpc10 <= 13'sd197/*197:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh3e] <= 8'h2;
                       end 
                      
                  13'sd197/*197:xpc10*/:  begin 
                       xpc10 <= 13'sd198/*198:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh3f] <= 8'h2;
                       end 
                      
                  13'sd198/*198:xpc10*/:  begin 
                       xpc10 <= 13'sd199/*199:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh40] <= 8'h1;
                       end 
                      
                  13'sd199/*199:xpc10*/:  begin 
                       xpc10 <= 13'sd200/*200:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh41] <= 8'h1;
                       end 
                      
                  13'sd200/*200:xpc10*/:  begin 
                       xpc10 <= 13'sd201/*201:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh42] <= 8'h1;
                       end 
                      
                  13'sd201/*201:xpc10*/:  begin 
                       xpc10 <= 13'sd202/*202:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh43] <= 8'h1;
                       end 
                      
                  13'sd202/*202:xpc10*/:  begin 
                       xpc10 <= 13'sd203/*203:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh44] <= 8'h1;
                       end 
                      
                  13'sd203/*203:xpc10*/:  begin 
                       xpc10 <= 13'sd204/*204:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh45] <= 8'h1;
                       end 
                      
                  13'sd204/*204:xpc10*/:  begin 
                       xpc10 <= 13'sd205/*205:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh46] <= 8'h1;
                       end 
                      
                  13'sd205/*205:xpc10*/:  begin 
                       xpc10 <= 13'sd206/*206:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh47] <= 8'h1;
                       end 
                      
                  13'sd206/*206:xpc10*/:  begin 
                       xpc10 <= 13'sd207/*207:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh48] <= 8'h1;
                       end 
                      
                  13'sd207/*207:xpc10*/:  begin 
                       xpc10 <= 13'sd208/*208:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh49] <= 8'h1;
                       end 
                      
                  13'sd208/*208:xpc10*/:  begin 
                       xpc10 <= 13'sd209/*209:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh4a] <= 8'h1;
                       end 
                      
                  13'sd209/*209:xpc10*/:  begin 
                       xpc10 <= 13'sd210/*210:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh4b] <= 8'h1;
                       end 
                      
                  13'sd210/*210:xpc10*/:  begin 
                       xpc10 <= 13'sd211/*211:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh4c] <= 8'h1;
                       end 
                      
                  13'sd211/*211:xpc10*/:  begin 
                       xpc10 <= 13'sd212/*212:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh4d] <= 8'h1;
                       end 
                      
                  13'sd212/*212:xpc10*/:  begin 
                       xpc10 <= 13'sd213/*213:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh4e] <= 8'h1;
                       end 
                      
                  13'sd213/*213:xpc10*/:  begin 
                       xpc10 <= 13'sd214/*214:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh4f] <= 8'h1;
                       end 
                      
                  13'sd214/*214:xpc10*/:  begin 
                       xpc10 <= 13'sd215/*215:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh50] <= 8'h1;
                       end 
                      
                  13'sd215/*215:xpc10*/:  begin 
                       xpc10 <= 13'sd216/*216:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh51] <= 8'h1;
                       end 
                      
                  13'sd216/*216:xpc10*/:  begin 
                       xpc10 <= 13'sd217/*217:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh52] <= 8'h1;
                       end 
                      
                  13'sd217/*217:xpc10*/:  begin 
                       xpc10 <= 13'sd218/*218:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh53] <= 8'h1;
                       end 
                      
                  13'sd218/*218:xpc10*/:  begin 
                       xpc10 <= 13'sd219/*219:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh54] <= 8'h1;
                       end 
                      
                  13'sd219/*219:xpc10*/:  begin 
                       xpc10 <= 13'sd220/*220:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh55] <= 8'h1;
                       end 
                      
                  13'sd220/*220:xpc10*/:  begin 
                       xpc10 <= 13'sd221/*221:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh56] <= 8'h1;
                       end 
                      
                  13'sd221/*221:xpc10*/:  begin 
                       xpc10 <= 13'sd222/*222:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh57] <= 8'h1;
                       end 
                      
                  13'sd222/*222:xpc10*/:  begin 
                       xpc10 <= 13'sd223/*223:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh58] <= 8'h1;
                       end 
                      
                  13'sd223/*223:xpc10*/:  begin 
                       xpc10 <= 13'sd224/*224:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh59] <= 8'h1;
                       end 
                      
                  13'sd224/*224:xpc10*/:  begin 
                       xpc10 <= 13'sd225/*225:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh5a] <= 8'h1;
                       end 
                      
                  13'sd225/*225:xpc10*/:  begin 
                       xpc10 <= 13'sd226/*226:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh5b] <= 8'h1;
                       end 
                      
                  13'sd226/*226:xpc10*/:  begin 
                       xpc10 <= 13'sd227/*227:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh5c] <= 8'h1;
                       end 
                      
                  13'sd227/*227:xpc10*/:  begin 
                       xpc10 <= 13'sd228/*228:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh5d] <= 8'h1;
                       end 
                      
                  13'sd228/*228:xpc10*/:  begin 
                       xpc10 <= 13'sd229/*229:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh5e] <= 8'h1;
                       end 
                      
                  13'sd229/*229:xpc10*/:  begin 
                       xpc10 <= 13'sd230/*230:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh5f] <= 8'h1;
                       end 
                      
                  13'sd230/*230:xpc10*/:  begin 
                       xpc10 <= 13'sd231/*231:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh60] <= 8'h1;
                       end 
                      
                  13'sd231/*231:xpc10*/:  begin 
                       xpc10 <= 13'sd232/*232:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh61] <= 8'h1;
                       end 
                      
                  13'sd232/*232:xpc10*/:  begin 
                       xpc10 <= 13'sd233/*233:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh62] <= 8'h1;
                       end 
                      
                  13'sd233/*233:xpc10*/:  begin 
                       xpc10 <= 13'sd234/*234:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh63] <= 8'h1;
                       end 
                      
                  13'sd234/*234:xpc10*/:  begin 
                       xpc10 <= 13'sd235/*235:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh64] <= 8'h1;
                       end 
                      
                  13'sd235/*235:xpc10*/:  begin 
                       xpc10 <= 13'sd236/*236:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh65] <= 8'h1;
                       end 
                      
                  13'sd236/*236:xpc10*/:  begin 
                       xpc10 <= 13'sd237/*237:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh66] <= 8'h1;
                       end 
                      
                  13'sd237/*237:xpc10*/:  begin 
                       xpc10 <= 13'sd238/*238:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh67] <= 8'h1;
                       end 
                      
                  13'sd238/*238:xpc10*/:  begin 
                       xpc10 <= 13'sd239/*239:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh68] <= 8'h1;
                       end 
                      
                  13'sd239/*239:xpc10*/:  begin 
                       xpc10 <= 13'sd240/*240:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh69] <= 8'h1;
                       end 
                      
                  13'sd240/*240:xpc10*/:  begin 
                       xpc10 <= 13'sd241/*241:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh6a] <= 8'h1;
                       end 
                      
                  13'sd241/*241:xpc10*/:  begin 
                       xpc10 <= 13'sd242/*242:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh6b] <= 8'h1;
                       end 
                      
                  13'sd242/*242:xpc10*/:  begin 
                       xpc10 <= 13'sd243/*243:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh6c] <= 8'h1;
                       end 
                      
                  13'sd243/*243:xpc10*/:  begin 
                       xpc10 <= 13'sd244/*244:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh6d] <= 8'h1;
                       end 
                      
                  13'sd244/*244:xpc10*/:  begin 
                       xpc10 <= 13'sd245/*245:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh6e] <= 8'h1;
                       end 
                      
                  13'sd245/*245:xpc10*/:  begin 
                       xpc10 <= 13'sd246/*246:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh6f] <= 8'h1;
                       end 
                      
                  13'sd246/*246:xpc10*/:  begin 
                       xpc10 <= 13'sd247/*247:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh70] <= 8'h1;
                       end 
                      
                  13'sd247/*247:xpc10*/:  begin 
                       xpc10 <= 13'sd248/*248:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh71] <= 8'h1;
                       end 
                      
                  13'sd248/*248:xpc10*/:  begin 
                       xpc10 <= 13'sd249/*249:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh72] <= 8'h1;
                       end 
                      
                  13'sd249/*249:xpc10*/:  begin 
                       xpc10 <= 13'sd250/*250:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh73] <= 8'h1;
                       end 
                      
                  13'sd250/*250:xpc10*/:  begin 
                       xpc10 <= 13'sd251/*251:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh74] <= 8'h1;
                       end 
                      
                  13'sd251/*251:xpc10*/:  begin 
                       xpc10 <= 13'sd252/*252:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh75] <= 8'h1;
                       end 
                      
                  13'sd252/*252:xpc10*/:  begin 
                       xpc10 <= 13'sd253/*253:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh76] <= 8'h1;
                       end 
                      
                  13'sd253/*253:xpc10*/:  begin 
                       xpc10 <= 13'sd254/*254:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh77] <= 8'h1;
                       end 
                      
                  13'sd254/*254:xpc10*/:  begin 
                       xpc10 <= 13'sd255/*255:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh78] <= 8'h1;
                       end 
                      
                  13'sd255/*255:xpc10*/:  begin 
                       xpc10 <= 13'sd256/*256:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh79] <= 8'h1;
                       end 
                      
                  13'sd256/*256:xpc10*/:  begin 
                       xpc10 <= 13'sd257/*257:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh7a] <= 8'h1;
                       end 
                      
                  13'sd257/*257:xpc10*/:  begin 
                       xpc10 <= 13'sd258/*258:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh7b] <= 8'h1;
                       end 
                      
                  13'sd258/*258:xpc10*/:  begin 
                       xpc10 <= 13'sd259/*259:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh7c] <= 8'h1;
                       end 
                      
                  13'sd259/*259:xpc10*/:  begin 
                       xpc10 <= 13'sd260/*260:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh7d] <= 8'h1;
                       end 
                      
                  13'sd260/*260:xpc10*/:  begin 
                       xpc10 <= 13'sd261/*261:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh7e] <= 8'h1;
                       end 
                      
                  13'sd261/*261:xpc10*/:  begin 
                       xpc10 <= 13'sd262/*262:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh7f] <= 8'h1;
                       end 
                      
                  13'sd262/*262:xpc10*/:  begin 
                       xpc10 <= 13'sd263/*263:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh80] <= 8'h0;
                       end 
                      
                  13'sd263/*263:xpc10*/:  begin 
                       xpc10 <= 13'sd264/*264:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh81] <= 8'h0;
                       end 
                      
                  13'sd264/*264:xpc10*/:  begin 
                       xpc10 <= 13'sd265/*265:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh82] <= 8'h0;
                       end 
                      
                  13'sd265/*265:xpc10*/:  begin 
                       xpc10 <= 13'sd266/*266:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh83] <= 8'h0;
                       end 
                      
                  13'sd266/*266:xpc10*/:  begin 
                       xpc10 <= 13'sd267/*267:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh84] <= 8'h0;
                       end 
                      
                  13'sd267/*267:xpc10*/:  begin 
                       xpc10 <= 13'sd268/*268:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh85] <= 8'h0;
                       end 
                      
                  13'sd268/*268:xpc10*/:  begin 
                       xpc10 <= 13'sd269/*269:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh86] <= 8'h0;
                       end 
                      
                  13'sd269/*269:xpc10*/:  begin 
                       xpc10 <= 13'sd270/*270:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh87] <= 8'h0;
                       end 
                      
                  13'sd270/*270:xpc10*/:  begin 
                       xpc10 <= 13'sd271/*271:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh88] <= 8'h0;
                       end 
                      
                  13'sd271/*271:xpc10*/:  begin 
                       xpc10 <= 13'sd272/*272:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh89] <= 8'h0;
                       end 
                      
                  13'sd272/*272:xpc10*/:  begin 
                       xpc10 <= 13'sd273/*273:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh8a] <= 8'h0;
                       end 
                      
                  13'sd273/*273:xpc10*/:  begin 
                       xpc10 <= 13'sd274/*274:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh8b] <= 8'h0;
                       end 
                      
                  13'sd274/*274:xpc10*/:  begin 
                       xpc10 <= 13'sd275/*275:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh8c] <= 8'h0;
                       end 
                      
                  13'sd275/*275:xpc10*/:  begin 
                       xpc10 <= 13'sd276/*276:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh8d] <= 8'h0;
                       end 
                      
                  13'sd276/*276:xpc10*/:  begin 
                       xpc10 <= 13'sd277/*277:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh8e] <= 8'h0;
                       end 
                      
                  13'sd277/*277:xpc10*/:  begin 
                       xpc10 <= 13'sd278/*278:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh8f] <= 8'h0;
                       end 
                      
                  13'sd278/*278:xpc10*/:  begin 
                       xpc10 <= 13'sd279/*279:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh90] <= 8'h0;
                       end 
                      
                  13'sd279/*279:xpc10*/:  begin 
                       xpc10 <= 13'sd280/*280:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh91] <= 8'h0;
                       end 
                      
                  13'sd280/*280:xpc10*/:  begin 
                       xpc10 <= 13'sd281/*281:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh92] <= 8'h0;
                       end 
                      
                  13'sd281/*281:xpc10*/:  begin 
                       xpc10 <= 13'sd282/*282:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh93] <= 8'h0;
                       end 
                      
                  13'sd282/*282:xpc10*/:  begin 
                       xpc10 <= 13'sd283/*283:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh94] <= 8'h0;
                       end 
                      
                  13'sd283/*283:xpc10*/:  begin 
                       xpc10 <= 13'sd284/*284:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh95] <= 8'h0;
                       end 
                      
                  13'sd284/*284:xpc10*/:  begin 
                       xpc10 <= 13'sd285/*285:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh96] <= 8'h0;
                       end 
                      
                  13'sd285/*285:xpc10*/:  begin 
                       xpc10 <= 13'sd286/*286:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh97] <= 8'h0;
                       end 
                      
                  13'sd286/*286:xpc10*/:  begin 
                       xpc10 <= 13'sd287/*287:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh98] <= 8'h0;
                       end 
                      
                  13'sd287/*287:xpc10*/:  begin 
                       xpc10 <= 13'sd288/*288:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh99] <= 8'h0;
                       end 
                      
                  13'sd288/*288:xpc10*/:  begin 
                       xpc10 <= 13'sd289/*289:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh9a] <= 8'h0;
                       end 
                      
                  13'sd289/*289:xpc10*/:  begin 
                       xpc10 <= 13'sd290/*290:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh9b] <= 8'h0;
                       end 
                      
                  13'sd290/*290:xpc10*/:  begin 
                       xpc10 <= 13'sd291/*291:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh9c] <= 8'h0;
                       end 
                      
                  13'sd291/*291:xpc10*/:  begin 
                       xpc10 <= 13'sd292/*292:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh9d] <= 8'h0;
                       end 
                      
                  13'sd292/*292:xpc10*/:  begin 
                       xpc10 <= 13'sd293/*293:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh9e] <= 8'h0;
                       end 
                      
                  13'sd293/*293:xpc10*/:  begin 
                       xpc10 <= 13'sd294/*294:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sh9f] <= 8'h0;
                       end 
                      
                  13'sd294/*294:xpc10*/:  begin 
                       xpc10 <= 13'sd295/*295:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sha0] <= 8'h0;
                       end 
                      
                  13'sd295/*295:xpc10*/:  begin 
                       xpc10 <= 13'sd296/*296:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sha1] <= 8'h0;
                       end 
                      
                  13'sd296/*296:xpc10*/:  begin 
                       xpc10 <= 13'sd297/*297:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sha2] <= 8'h0;
                       end 
                      
                  13'sd297/*297:xpc10*/:  begin 
                       xpc10 <= 13'sd298/*298:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sha3] <= 8'h0;
                       end 
                      
                  13'sd298/*298:xpc10*/:  begin 
                       xpc10 <= 13'sd299/*299:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sha4] <= 8'h0;
                       end 
                      
                  13'sd299/*299:xpc10*/:  begin 
                       xpc10 <= 13'sd300/*300:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sha5] <= 8'h0;
                       end 
                      
                  13'sd300/*300:xpc10*/:  begin 
                       xpc10 <= 13'sd301/*301:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sha6] <= 8'h0;
                       end 
                      
                  13'sd301/*301:xpc10*/:  begin 
                       xpc10 <= 13'sd302/*302:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sha7] <= 8'h0;
                       end 
                      
                  13'sd302/*302:xpc10*/:  begin 
                       xpc10 <= 13'sd303/*303:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sha8] <= 8'h0;
                       end 
                      
                  13'sd303/*303:xpc10*/:  begin 
                       xpc10 <= 13'sd304/*304:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sha9] <= 8'h0;
                       end 
                      
                  13'sd304/*304:xpc10*/:  begin 
                       xpc10 <= 13'sd305/*305:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shaa] <= 8'h0;
                       end 
                      
                  13'sd305/*305:xpc10*/:  begin 
                       xpc10 <= 13'sd306/*306:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shab] <= 8'h0;
                       end 
                      
                  13'sd306/*306:xpc10*/:  begin 
                       xpc10 <= 13'sd307/*307:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shac] <= 8'h0;
                       end 
                      
                  13'sd307/*307:xpc10*/:  begin 
                       xpc10 <= 13'sd308/*308:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shad] <= 8'h0;
                       end 
                      
                  13'sd308/*308:xpc10*/:  begin 
                       xpc10 <= 13'sd309/*309:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shae] <= 8'h0;
                       end 
                      
                  13'sd309/*309:xpc10*/:  begin 
                       xpc10 <= 13'sd310/*310:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shaf] <= 8'h0;
                       end 
                      
                  13'sd310/*310:xpc10*/:  begin 
                       xpc10 <= 13'sd311/*311:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shb0] <= 8'h0;
                       end 
                      
                  13'sd311/*311:xpc10*/:  begin 
                       xpc10 <= 13'sd312/*312:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shb1] <= 8'h0;
                       end 
                      
                  13'sd312/*312:xpc10*/:  begin 
                       xpc10 <= 13'sd313/*313:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shb2] <= 8'h0;
                       end 
                      
                  13'sd313/*313:xpc10*/:  begin 
                       xpc10 <= 13'sd314/*314:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shb3] <= 8'h0;
                       end 
                      
                  13'sd314/*314:xpc10*/:  begin 
                       xpc10 <= 13'sd315/*315:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shb4] <= 8'h0;
                       end 
                      
                  13'sd315/*315:xpc10*/:  begin 
                       xpc10 <= 13'sd316/*316:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shb5] <= 8'h0;
                       end 
                      
                  13'sd316/*316:xpc10*/:  begin 
                       xpc10 <= 13'sd317/*317:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shb6] <= 8'h0;
                       end 
                      
                  13'sd317/*317:xpc10*/:  begin 
                       xpc10 <= 13'sd318/*318:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shb7] <= 8'h0;
                       end 
                      
                  13'sd318/*318:xpc10*/:  begin 
                       xpc10 <= 13'sd319/*319:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shb8] <= 8'h0;
                       end 
                      
                  13'sd319/*319:xpc10*/:  begin 
                       xpc10 <= 13'sd320/*320:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shb9] <= 8'h0;
                       end 
                      
                  13'sd320/*320:xpc10*/:  begin 
                       xpc10 <= 13'sd321/*321:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shba] <= 8'h0;
                       end 
                      
                  13'sd321/*321:xpc10*/:  begin 
                       xpc10 <= 13'sd322/*322:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shbb] <= 8'h0;
                       end 
                      
                  13'sd322/*322:xpc10*/:  begin 
                       xpc10 <= 13'sd323/*323:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shbc] <= 8'h0;
                       end 
                      
                  13'sd323/*323:xpc10*/:  begin 
                       xpc10 <= 13'sd324/*324:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shbd] <= 8'h0;
                       end 
                      
                  13'sd324/*324:xpc10*/:  begin 
                       xpc10 <= 13'sd325/*325:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shbe] <= 8'h0;
                       end 
                      
                  13'sd325/*325:xpc10*/:  begin 
                       xpc10 <= 13'sd326/*326:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shbf] <= 8'h0;
                       end 
                      
                  13'sd326/*326:xpc10*/:  begin 
                       xpc10 <= 13'sd327/*327:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shc0] <= 8'h0;
                       end 
                      
                  13'sd327/*327:xpc10*/:  begin 
                       xpc10 <= 13'sd328/*328:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shc1] <= 8'h0;
                       end 
                      
                  13'sd328/*328:xpc10*/:  begin 
                       xpc10 <= 13'sd329/*329:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shc2] <= 8'h0;
                       end 
                      
                  13'sd329/*329:xpc10*/:  begin 
                       xpc10 <= 13'sd330/*330:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shc3] <= 8'h0;
                       end 
                      
                  13'sd330/*330:xpc10*/:  begin 
                       xpc10 <= 13'sd331/*331:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shc4] <= 8'h0;
                       end 
                      
                  13'sd331/*331:xpc10*/:  begin 
                       xpc10 <= 13'sd332/*332:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shc5] <= 8'h0;
                       end 
                      
                  13'sd332/*332:xpc10*/:  begin 
                       xpc10 <= 13'sd333/*333:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shc6] <= 8'h0;
                       end 
                      
                  13'sd333/*333:xpc10*/:  begin 
                       xpc10 <= 13'sd334/*334:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shc7] <= 8'h0;
                       end 
                      
                  13'sd334/*334:xpc10*/:  begin 
                       xpc10 <= 13'sd335/*335:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shc8] <= 8'h0;
                       end 
                      
                  13'sd335/*335:xpc10*/:  begin 
                       xpc10 <= 13'sd336/*336:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shc9] <= 8'h0;
                       end 
                      
                  13'sd336/*336:xpc10*/:  begin 
                       xpc10 <= 13'sd337/*337:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shca] <= 8'h0;
                       end 
                      
                  13'sd337/*337:xpc10*/:  begin 
                       xpc10 <= 13'sd338/*338:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shcb] <= 8'h0;
                       end 
                      
                  13'sd338/*338:xpc10*/:  begin 
                       xpc10 <= 13'sd339/*339:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shcc] <= 8'h0;
                       end 
                      
                  13'sd339/*339:xpc10*/:  begin 
                       xpc10 <= 13'sd340/*340:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shcd] <= 8'h0;
                       end 
                      
                  13'sd340/*340:xpc10*/:  begin 
                       xpc10 <= 13'sd341/*341:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shce] <= 8'h0;
                       end 
                      
                  13'sd341/*341:xpc10*/:  begin 
                       xpc10 <= 13'sd342/*342:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shcf] <= 8'h0;
                       end 
                      
                  13'sd342/*342:xpc10*/:  begin 
                       xpc10 <= 13'sd343/*343:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shd0] <= 8'h0;
                       end 
                      
                  13'sd343/*343:xpc10*/:  begin 
                       xpc10 <= 13'sd344/*344:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shd1] <= 8'h0;
                       end 
                      
                  13'sd344/*344:xpc10*/:  begin 
                       xpc10 <= 13'sd345/*345:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shd2] <= 8'h0;
                       end 
                      
                  13'sd345/*345:xpc10*/:  begin 
                       xpc10 <= 13'sd346/*346:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shd3] <= 8'h0;
                       end 
                      
                  13'sd346/*346:xpc10*/:  begin 
                       xpc10 <= 13'sd347/*347:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shd4] <= 8'h0;
                       end 
                      
                  13'sd347/*347:xpc10*/:  begin 
                       xpc10 <= 13'sd348/*348:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shd5] <= 8'h0;
                       end 
                      
                  13'sd348/*348:xpc10*/:  begin 
                       xpc10 <= 13'sd349/*349:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shd6] <= 8'h0;
                       end 
                      
                  13'sd349/*349:xpc10*/:  begin 
                       xpc10 <= 13'sd350/*350:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shd7] <= 8'h0;
                       end 
                      
                  13'sd350/*350:xpc10*/:  begin 
                       xpc10 <= 13'sd351/*351:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shd8] <= 8'h0;
                       end 
                      
                  13'sd351/*351:xpc10*/:  begin 
                       xpc10 <= 13'sd352/*352:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shd9] <= 8'h0;
                       end 
                      
                  13'sd352/*352:xpc10*/:  begin 
                       xpc10 <= 13'sd353/*353:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shda] <= 8'h0;
                       end 
                      
                  13'sd353/*353:xpc10*/:  begin 
                       xpc10 <= 13'sd354/*354:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shdb] <= 8'h0;
                       end 
                      
                  13'sd354/*354:xpc10*/:  begin 
                       xpc10 <= 13'sd355/*355:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shdc] <= 8'h0;
                       end 
                      
                  13'sd355/*355:xpc10*/:  begin 
                       xpc10 <= 13'sd356/*356:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shdd] <= 8'h0;
                       end 
                      
                  13'sd356/*356:xpc10*/:  begin 
                       xpc10 <= 13'sd357/*357:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shde] <= 8'h0;
                       end 
                      
                  13'sd357/*357:xpc10*/:  begin 
                       xpc10 <= 13'sd358/*358:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shdf] <= 8'h0;
                       end 
                      
                  13'sd358/*358:xpc10*/:  begin 
                       xpc10 <= 13'sd359/*359:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'she0] <= 8'h0;
                       end 
                      
                  13'sd359/*359:xpc10*/:  begin 
                       xpc10 <= 13'sd360/*360:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'she1] <= 8'h0;
                       end 
                      
                  13'sd360/*360:xpc10*/:  begin 
                       xpc10 <= 13'sd361/*361:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'she2] <= 8'h0;
                       end 
                      
                  13'sd361/*361:xpc10*/:  begin 
                       xpc10 <= 13'sd362/*362:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'she3] <= 8'h0;
                       end 
                      
                  13'sd362/*362:xpc10*/:  begin 
                       xpc10 <= 13'sd363/*363:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'she4] <= 8'h0;
                       end 
                      
                  13'sd363/*363:xpc10*/:  begin 
                       xpc10 <= 13'sd364/*364:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'she5] <= 8'h0;
                       end 
                      
                  13'sd364/*364:xpc10*/:  begin 
                       xpc10 <= 13'sd365/*365:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'she6] <= 8'h0;
                       end 
                      
                  13'sd365/*365:xpc10*/:  begin 
                       xpc10 <= 13'sd366/*366:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'she7] <= 8'h0;
                       end 
                      
                  13'sd366/*366:xpc10*/:  begin 
                       xpc10 <= 13'sd367/*367:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'she8] <= 8'h0;
                       end 
                      
                  13'sd367/*367:xpc10*/:  begin 
                       xpc10 <= 13'sd368/*368:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'she9] <= 8'h0;
                       end 
                      
                  13'sd368/*368:xpc10*/:  begin 
                       xpc10 <= 13'sd369/*369:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shea] <= 8'h0;
                       end 
                      
                  13'sd369/*369:xpc10*/:  begin 
                       xpc10 <= 13'sd370/*370:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'sheb] <= 8'h0;
                       end 
                      
                  13'sd370/*370:xpc10*/:  begin 
                       xpc10 <= 13'sd371/*371:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shec] <= 8'h0;
                       end 
                      
                  13'sd371/*371:xpc10*/:  begin 
                       xpc10 <= 13'sd372/*372:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shed] <= 8'h0;
                       end 
                      
                  13'sd372/*372:xpc10*/:  begin 
                       xpc10 <= 13'sd373/*373:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shee] <= 8'h0;
                       end 
                      
                  13'sd373/*373:xpc10*/:  begin 
                       xpc10 <= 13'sd374/*374:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shef] <= 8'h0;
                       end 
                      
                  13'sd374/*374:xpc10*/:  begin 
                       xpc10 <= 13'sd375/*375:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shf0] <= 8'h0;
                       end 
                      
                  13'sd375/*375:xpc10*/:  begin 
                       xpc10 <= 13'sd376/*376:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shf1] <= 8'h0;
                       end 
                      
                  13'sd376/*376:xpc10*/:  begin 
                       xpc10 <= 13'sd377/*377:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shf2] <= 8'h0;
                       end 
                      
                  13'sd377/*377:xpc10*/:  begin 
                       xpc10 <= 13'sd378/*378:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shf3] <= 8'h0;
                       end 
                      
                  13'sd378/*378:xpc10*/:  begin 
                       xpc10 <= 13'sd379/*379:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shf4] <= 8'h0;
                       end 
                      
                  13'sd379/*379:xpc10*/:  begin 
                       xpc10 <= 13'sd380/*380:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shf5] <= 8'h0;
                       end 
                      
                  13'sd380/*380:xpc10*/:  begin 
                       xpc10 <= 13'sd381/*381:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shf6] <= 8'h0;
                       end 
                      
                  13'sd381/*381:xpc10*/:  begin 
                       xpc10 <= 13'sd382/*382:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shf7] <= 8'h0;
                       end 
                      
                  13'sd382/*382:xpc10*/:  begin 
                       xpc10 <= 13'sd383/*383:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shf8] <= 8'h0;
                       end 
                      
                  13'sd383/*383:xpc10*/:  begin 
                       xpc10 <= 13'sd384/*384:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shf9] <= 8'h0;
                       end 
                      
                  13'sd384/*384:xpc10*/:  begin 
                       xpc10 <= 13'sd385/*385:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shfa] <= 8'h0;
                       end 
                      
                  13'sd385/*385:xpc10*/:  begin 
                       xpc10 <= 13'sd386/*386:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shfb] <= 8'h0;
                       end 
                      
                  13'sd386/*386:xpc10*/:  begin 
                       xpc10 <= 13'sd387/*387:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shfc] <= 8'h0;
                       end 
                      
                  13'sd387/*387:xpc10*/:  begin 
                       xpc10 <= 13'sd388/*388:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shfd] <= 8'h0;
                       end 
                      
                  13'sd388/*388:xpc10*/:  begin 
                       xpc10 <= 13'sd389/*389:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shfe] <= 8'h0;
                       end 
                      
                  13'sd389/*389:xpc10*/:  begin 
                       xpc10 <= 13'sd390/*390:xpc10*/;
                       A_8_US_CC_SCALbx16_ARA0[64'shff] <= 8'h0;
                       end 
                      
                  13'sd415/*415:xpc10*/:  xpc10 <= 13'sd416/*416:xpc10*/;

                  13'sd417/*417:xpc10*/:  begin 
                       xpc10 <= 13'sd418/*418:xpc10*/;
                       Tdbm0_3_V_0 <= 32'sd0;
                       end 
                      
                  13'sd418/*418:xpc10*/:  begin 
                       xpc10 <= 13'sd419/*419:xpc10*/;
                       Tdbm0_3_V_1 <= 32'sd1;
                       end 
                      
                  13'sd426/*426:xpc10*/:  begin 
                       xpc10 <= 13'sd427/*427:xpc10*/;
                       Tdsi1_5_V_0 <= $unsigned(A_64_US_CC_SCALbx12_ARB0[Tdbm0_3_V_1]);
                       end 
                      
                  13'sd427/*427:xpc10*/:  begin 
                       xpc10 <= 13'sd428/*428:xpc10*/;
                       Tdsi1_5_V_1 <= $unsigned(A_64_US_CC_SCALbx12_ARB0[Tdbm0_3_V_1]);
                       end 
                      
                  13'sd428/*428:xpc10*/:  begin 
                       xpc10 <= 13'sd429/*429:xpc10*/;
                       Tdsi1_5_V_2 <= 32'sd1;
                       end 
                      
                  13'sd429/*429:xpc10*/:  begin 
                       xpc10 <= 13'sd430/*430:xpc10*/;
                       Tsfl0_9_V_8 <= 64'h0;
                       end 
                      
                  13'sd430/*430:xpc10*/:  begin 
                       xpc10 <= 13'sd431/*431:xpc10*/;
                       Tsfl0_9_V_9 <= 64'h0;
                       end 
                      
                  13'sd431/*431:xpc10*/:  begin 
                       xpc10 <= 13'sd432/*432:xpc10*/;
                       Tsfl0_9_V_6 <= 64'shf_ffff_ffff_ffff&A_64_US_CC_SCALbx12_ARB0[Tdbm0_3_V_1];
                       end 
                      
                  13'sd432/*432:xpc10*/:  begin 
                       xpc10 <= 13'sd433/*433:xpc10*/;
                       Tsfl0_9_V_3 <= rtl_signed_bitextract2(64'sh7ff&(A_64_US_CC_SCALbx12_ARB0[Tdbm0_3_V_1]>>32'sd52));
                       end 
                      
                  13'sd437/*437:xpc10*/:  begin 
                       xpc10 <= 13'sd438/*438:xpc10*/;
                       Tse0_SPILL_256 <= 32'sd1;
                       end 
                      
                  13'sd441/*441:xpc10*/:  begin 
                       xpc10 <= 13'sd442/*442:xpc10*/;
                       Tsfl0_9_V_0 <= rtl_unsigned_bitextract4(Tse0_SPILL_256);
                       end 
                      
                  13'sd442/*442:xpc10*/:  begin 
                       xpc10 <= 13'sd443/*443:xpc10*/;
                       Tsfl0_9_V_7 <= 64'shf_ffff_ffff_ffff&A_64_US_CC_SCALbx12_ARB0[Tdbm0_3_V_1];
                       end 
                      
                  13'sd443/*443:xpc10*/:  begin 
                       xpc10 <= 13'sd444/*444:xpc10*/;
                       Tsfl0_9_V_4 <= rtl_signed_bitextract2(64'sh7ff&(A_64_US_CC_SCALbx12_ARB0[Tdbm0_3_V_1]>>32'sd52));
                       end 
                      
                  13'sd448/*448:xpc10*/:  begin 
                       xpc10 <= 13'sd449/*449:xpc10*/;
                       Tse0SPILL10_256 <= 32'sd1;
                       end 
                      
                  13'sd452/*452:xpc10*/:  begin 
                       xpc10 <= 13'sd453/*453:xpc10*/;
                       Tsfl0_9_V_1 <= rtl_unsigned_bitextract4(Tse0SPILL10_256);
                       end 
                      
                  13'sd453/*453:xpc10*/:  begin 
                       xpc10 <= 13'sd454/*454:xpc10*/;
                       Tsfl0_9_V_2 <= rtl_unsigned_bitextract12(Tsfl0_9_V_0^Tsfl0_9_V_1);
                       end 
                      endcase
              if ((13'sd0/*0:xpc10*/==xpc10))  xpc10 <= 13'sd1/*1:xpc10*/;
                  if ((13'sd1/*1:xpc10*/==xpc10))  xpc10 <= 13'sd2/*2:xpc10*/;
                  if ((13'sd2/*2:xpc10*/==xpc10))  xpc10 <= 13'sd3/*3:xpc10*/;
                  if ((13'sd3/*3:xpc10*/==xpc10))  xpc10 <= 13'sd4/*4:xpc10*/;
                  if ((13'sd4/*4:xpc10*/==xpc10))  xpc10 <= 13'sd5/*5:xpc10*/;
                  if ((13'sd5/*5:xpc10*/==xpc10))  xpc10 <= 13'sd6/*6:xpc10*/;
                  if ((13'sd6/*6:xpc10*/==xpc10))  xpc10 <= 13'sd7/*7:xpc10*/;
                  if ((13'sd7/*7:xpc10*/==xpc10))  xpc10 <= 13'sd8/*8:xpc10*/;
                  if ((13'sd8/*8:xpc10*/==xpc10))  xpc10 <= 13'sd9/*9:xpc10*/;
                  if ((13'sd9/*9:xpc10*/==xpc10))  xpc10 <= 13'sd10/*10:xpc10*/;
                  if ((13'sd10/*10:xpc10*/==xpc10))  xpc10 <= 13'sd11/*11:xpc10*/;
                  if ((13'sd11/*11:xpc10*/==xpc10))  xpc10 <= 13'sd12/*12:xpc10*/;
                  if ((13'sd12/*12:xpc10*/==xpc10))  xpc10 <= 13'sd13/*13:xpc10*/;
                  if ((13'sd13/*13:xpc10*/==xpc10))  xpc10 <= 13'sd14/*14:xpc10*/;
                  if ((13'sd14/*14:xpc10*/==xpc10))  xpc10 <= 13'sd15/*15:xpc10*/;
                  if ((13'sd15/*15:xpc10*/==xpc10))  xpc10 <= 13'sd16/*16:xpc10*/;
                  if ((13'sd16/*16:xpc10*/==xpc10))  xpc10 <= 13'sd17/*17:xpc10*/;
                  if ((13'sd17/*17:xpc10*/==xpc10))  xpc10 <= 13'sd18/*18:xpc10*/;
                  if ((13'sd18/*18:xpc10*/==xpc10))  xpc10 <= 13'sd19/*19:xpc10*/;
                  if ((13'sd19/*19:xpc10*/==xpc10))  xpc10 <= 13'sd20/*20:xpc10*/;
                  if ((13'sd20/*20:xpc10*/==xpc10))  xpc10 <= 13'sd21/*21:xpc10*/;
                  if ((13'sd21/*21:xpc10*/==xpc10))  xpc10 <= 13'sd22/*22:xpc10*/;
                  if ((13'sd22/*22:xpc10*/==xpc10))  xpc10 <= 13'sd23/*23:xpc10*/;
                  if ((13'sd23/*23:xpc10*/==xpc10))  xpc10 <= 13'sd24/*24:xpc10*/;
                  if ((13'sd24/*24:xpc10*/==xpc10))  xpc10 <= 13'sd25/*25:xpc10*/;
                  if ((13'sd25/*25:xpc10*/==xpc10))  xpc10 <= 13'sd26/*26:xpc10*/;
                  if ((13'sd26/*26:xpc10*/==xpc10))  xpc10 <= 13'sd27/*27:xpc10*/;
                  if ((13'sd27/*27:xpc10*/==xpc10))  xpc10 <= 13'sd28/*28:xpc10*/;
                  if ((13'sd28/*28:xpc10*/==xpc10))  xpc10 <= 13'sd29/*29:xpc10*/;
                  if ((13'sd29/*29:xpc10*/==xpc10))  xpc10 <= 13'sd30/*30:xpc10*/;
                  if ((13'sd30/*30:xpc10*/==xpc10))  xpc10 <= 13'sd31/*31:xpc10*/;
                  if ((13'sd31/*31:xpc10*/==xpc10))  xpc10 <= 13'sd32/*32:xpc10*/;
                  if ((13'sd32/*32:xpc10*/==xpc10))  xpc10 <= 13'sd33/*33:xpc10*/;
                  if ((13'sd33/*33:xpc10*/==xpc10))  xpc10 <= 13'sd34/*34:xpc10*/;
                  if ((13'sd34/*34:xpc10*/==xpc10))  xpc10 <= 13'sd35/*35:xpc10*/;
                  if ((13'sd35/*35:xpc10*/==xpc10))  xpc10 <= 13'sd36/*36:xpc10*/;
                  if ((13'sd36/*36:xpc10*/==xpc10))  xpc10 <= 13'sd37/*37:xpc10*/;
                  if ((13'sd37/*37:xpc10*/==xpc10))  xpc10 <= 13'sd38/*38:xpc10*/;
                  if ((13'sd38/*38:xpc10*/==xpc10))  xpc10 <= 13'sd39/*39:xpc10*/;
                  if ((13'sd39/*39:xpc10*/==xpc10))  xpc10 <= 13'sd40/*40:xpc10*/;
                  if ((13'sd40/*40:xpc10*/==xpc10))  xpc10 <= 13'sd41/*41:xpc10*/;
                  if ((13'sd41/*41:xpc10*/==xpc10))  xpc10 <= 13'sd42/*42:xpc10*/;
                  if ((13'sd42/*42:xpc10*/==xpc10))  xpc10 <= 13'sd43/*43:xpc10*/;
                  if ((13'sd43/*43:xpc10*/==xpc10))  xpc10 <= 13'sd44/*44:xpc10*/;
                  if ((13'sd44/*44:xpc10*/==xpc10))  xpc10 <= 13'sd45/*45:xpc10*/;
                  if ((13'sd45/*45:xpc10*/==xpc10))  xpc10 <= 13'sd46/*46:xpc10*/;
                  if ((13'sd82/*82:xpc10*/==xpc10))  xpc10 <= 13'sd83/*83:xpc10*/;
                  if ((13'sd83/*83:xpc10*/==xpc10))  xpc10 <= 13'sd84/*84:xpc10*/;
                  if ((13'sd84/*84:xpc10*/==xpc10))  xpc10 <= 13'sd85/*85:xpc10*/;
                  if ((13'sd121/*121:xpc10*/==xpc10))  xpc10 <= 13'sd122/*122:xpc10*/;
                  if ((13'sd123/*123:xpc10*/==xpc10))  xpc10 <= 13'sd124/*124:xpc10*/;
                  if ((13'sd124/*124:xpc10*/==xpc10))  xpc10 <= 13'sd125/*125:xpc10*/;
                  if ((13'sd125/*125:xpc10*/==xpc10))  xpc10 <= 13'sd126/*126:xpc10*/;
                  if ((13'sd126/*126:xpc10*/==xpc10))  xpc10 <= 13'sd127/*127:xpc10*/;
                  if ((13'sd127/*127:xpc10*/==xpc10))  xpc10 <= 13'sd128/*128:xpc10*/;
                  if ((13'sd128/*128:xpc10*/==xpc10))  xpc10 <= 13'sd129/*129:xpc10*/;
                  if ((13'sd129/*129:xpc10*/==xpc10))  xpc10 <= 13'sd130/*130:xpc10*/;
                  if ((13'sd130/*130:xpc10*/==xpc10))  xpc10 <= 13'sd131/*131:xpc10*/;
                  if ((13'sd131/*131:xpc10*/==xpc10))  xpc10 <= 13'sd132/*132:xpc10*/;
                  if ((13'sd132/*132:xpc10*/==xpc10))  xpc10 <= 13'sd133/*133:xpc10*/;
                  if ((13'sd133/*133:xpc10*/==xpc10))  xpc10 <= 13'sd134/*134:xpc10*/;
                  if ((13'sd390/*390:xpc10*/==xpc10))  xpc10 <= 13'sd391/*391:xpc10*/;
                  if ((13'sd391/*391:xpc10*/==xpc10))  xpc10 <= 13'sd392/*392:xpc10*/;
                  if ((13'sd392/*392:xpc10*/==xpc10))  xpc10 <= 13'sd393/*393:xpc10*/;
                  if ((13'sd393/*393:xpc10*/==xpc10))  xpc10 <= 13'sd394/*394:xpc10*/;
                  if ((13'sd394/*394:xpc10*/==xpc10))  xpc10 <= 13'sd395/*395:xpc10*/;
                  if ((13'sd395/*395:xpc10*/==xpc10))  xpc10 <= 13'sd396/*396:xpc10*/;
                  if ((13'sd396/*396:xpc10*/==xpc10))  xpc10 <= 13'sd397/*397:xpc10*/;
                  if ((13'sd397/*397:xpc10*/==xpc10))  xpc10 <= 13'sd398/*398:xpc10*/;
                  if ((13'sd398/*398:xpc10*/==xpc10))  xpc10 <= 13'sd399/*399:xpc10*/;
                  if ((13'sd399/*399:xpc10*/==xpc10))  xpc10 <= 13'sd400/*400:xpc10*/;
                  if ((13'sd400/*400:xpc10*/==xpc10))  xpc10 <= 13'sd401/*401:xpc10*/;
                  if ((13'sd401/*401:xpc10*/==xpc10))  xpc10 <= 13'sd402/*402:xpc10*/;
                  if ((13'sd402/*402:xpc10*/==xpc10))  xpc10 <= 13'sd403/*403:xpc10*/;
                  if ((13'sd403/*403:xpc10*/==xpc10))  xpc10 <= 13'sd404/*404:xpc10*/;
                  if ((13'sd404/*404:xpc10*/==xpc10))  xpc10 <= 13'sd405/*405:xpc10*/;
                  if ((13'sd405/*405:xpc10*/==xpc10))  xpc10 <= 13'sd406/*406:xpc10*/;
                  if ((13'sd406/*406:xpc10*/==xpc10))  xpc10 <= 13'sd407/*407:xpc10*/;
                  if ((13'sd407/*407:xpc10*/==xpc10))  xpc10 <= 13'sd408/*408:xpc10*/;
                  if ((13'sd408/*408:xpc10*/==xpc10))  xpc10 <= 13'sd409/*409:xpc10*/;
                  if ((13'sd409/*409:xpc10*/==xpc10))  xpc10 <= 13'sd410/*410:xpc10*/;
                  if ((13'sd410/*410:xpc10*/==xpc10))  xpc10 <= 13'sd411/*411:xpc10*/;
                  if ((13'sd411/*411:xpc10*/==xpc10))  xpc10 <= 13'sd412/*412:xpc10*/;
                  if ((13'sd412/*412:xpc10*/==xpc10))  xpc10 <= 13'sd413/*413:xpc10*/;
                  if ((13'sd413/*413:xpc10*/==xpc10))  xpc10 <= 13'sd414/*414:xpc10*/;
                  if ((13'sd414/*414:xpc10*/==xpc10))  xpc10 <= 13'sd415/*415:xpc10*/;
                  if ((13'sd416/*416:xpc10*/==xpc10))  xpc10 <= 13'sd417/*417:xpc10*/;
                  if ((13'sd419/*419:xpc10*/==xpc10))  xpc10 <= 13'sd420/*420:xpc10*/;
                  if ((13'sd420/*420:xpc10*/==xpc10))  xpc10 <= 13'sd421/*421:xpc10*/;
                  if ((13'sd421/*421:xpc10*/==xpc10))  xpc10 <= 13'sd422/*422:xpc10*/;
                  if ((13'sd422/*422:xpc10*/==xpc10))  xpc10 <= 13'sd423/*423:xpc10*/;
                  if ((13'sd423/*423:xpc10*/==xpc10))  xpc10 <= 13'sd424/*424:xpc10*/;
                  if ((13'sd424/*424:xpc10*/==xpc10))  xpc10 <= 13'sd425/*425:xpc10*/;
                  if ((13'sd425/*425:xpc10*/==xpc10))  xpc10 <= 13'sd426/*426:xpc10*/;
                  if ((13'sd434/*434:xpc10*/==xpc10))  xpc10 <= 13'sd435/*435:xpc10*/;
                  if ((13'sd435/*435:xpc10*/==xpc10))  xpc10 <= 13'sd436/*436:xpc10*/;
                  if ((13'sd436/*436:xpc10*/==xpc10))  xpc10 <= 13'sd437/*437:xpc10*/;
                  if ((13'sd438/*438:xpc10*/==xpc10))  xpc10 <= 13'sd439/*439:xpc10*/;
                  if ((13'sd439/*439:xpc10*/==xpc10))  xpc10 <= 13'sd440/*440:xpc10*/;
                  if ((13'sd440/*440:xpc10*/==xpc10))  xpc10 <= 13'sd441/*441:xpc10*/;
                  if ((13'sd445/*445:xpc10*/==xpc10))  xpc10 <= 13'sd446/*446:xpc10*/;
                  if ((13'sd446/*446:xpc10*/==xpc10))  xpc10 <= 13'sd447/*447:xpc10*/;
                  if ((13'sd447/*447:xpc10*/==xpc10))  xpc10 <= 13'sd448/*448:xpc10*/;
                  if ((13'sd449/*449:xpc10*/==xpc10))  xpc10 <= 13'sd450/*450:xpc10*/;
                  if ((13'sd450/*450:xpc10*/==xpc10))  xpc10 <= 13'sd451/*451:xpc10*/;
                  if ((13'sd451/*451:xpc10*/==xpc10))  xpc10 <= 13'sd452/*452:xpc10*/;
                  if ((13'sd455/*455:xpc10*/==xpc10))  xpc10 <= 13'sd456/*456:xpc10*/;
                  if ((13'sd456/*456:xpc10*/==xpc10))  xpc10 <= 13'sd457/*457:xpc10*/;
                  if ((13'sd457/*457:xpc10*/==xpc10))  xpc10 <= 13'sd458/*458:xpc10*/;
                  if ((13'sd459/*459:xpc10*/==xpc10))  xpc10 <= 13'sd460/*460:xpc10*/;
                  if ((13'sd460/*460:xpc10*/==xpc10))  xpc10 <= 13'sd461/*461:xpc10*/;
                  if ((13'sd461/*461:xpc10*/==xpc10))  xpc10 <= 13'sd462/*462:xpc10*/;
                  if ((13'sd463/*463:xpc10*/==xpc10))  xpc10 <= 13'sd464/*464:xpc10*/;
                  if ((13'sd464/*464:xpc10*/==xpc10))  xpc10 <= 13'sd465/*465:xpc10*/;
                  if ((13'sd465/*465:xpc10*/==xpc10))  xpc10 <= 13'sd466/*466:xpc10*/;
                  if ((13'sd467/*467:xpc10*/==xpc10))  xpc10 <= 13'sd468/*468:xpc10*/;
                  if ((13'sd468/*468:xpc10*/==xpc10))  xpc10 <= 13'sd469/*469:xpc10*/;
                  if ((13'sd469/*469:xpc10*/==xpc10))  xpc10 <= 13'sd470/*470:xpc10*/;
                  if ((13'sd473/*473:xpc10*/==xpc10))  xpc10 <= 13'sd474/*474:xpc10*/;
                  if ((13'sd474/*474:xpc10*/==xpc10))  xpc10 <= 13'sd475/*475:xpc10*/;
                  if ((13'sd475/*475:xpc10*/==xpc10))  xpc10 <= 13'sd476/*476:xpc10*/;
                  if ((13'sd477/*477:xpc10*/==xpc10))  xpc10 <= 13'sd478/*478:xpc10*/;
                  if ((13'sd478/*478:xpc10*/==xpc10))  xpc10 <= 13'sd479/*479:xpc10*/;
                  if ((13'sd479/*479:xpc10*/==xpc10))  xpc10 <= 13'sd480/*480:xpc10*/;
                  if ((13'sd483/*483:xpc10*/==xpc10))  xpc10 <= 13'sd484/*484:xpc10*/;
                  if ((13'sd484/*484:xpc10*/==xpc10))  xpc10 <= 13'sd485/*485:xpc10*/;
                  if ((13'sd485/*485:xpc10*/==xpc10))  xpc10 <= 13'sd486/*486:xpc10*/;
                  if ((13'sd487/*487:xpc10*/==xpc10))  xpc10 <= 13'sd488/*488:xpc10*/;
                  if ((13'sd488/*488:xpc10*/==xpc10))  xpc10 <= 13'sd489/*489:xpc10*/;
                  if ((13'sd489/*489:xpc10*/==xpc10))  xpc10 <= 13'sd490/*490:xpc10*/;
                  if ((13'sd494/*494:xpc10*/==xpc10))  xpc10 <= 13'sd495/*495:xpc10*/;
                  if ((13'sd495/*495:xpc10*/==xpc10))  xpc10 <= 13'sd496/*496:xpc10*/;
                  if ((13'sd496/*496:xpc10*/==xpc10))  xpc10 <= 13'sd497/*497:xpc10*/;
                  if ((13'sd497/*497:xpc10*/==xpc10))  xpc10 <= 13'sd498/*498:xpc10*/;
                  if ((13'sd498/*498:xpc10*/==xpc10))  xpc10 <= 13'sd499/*499:xpc10*/;
                  if ((13'sd499/*499:xpc10*/==xpc10))  xpc10 <= 13'sd500/*500:xpc10*/;
                  if ((13'sd500/*500:xpc10*/==xpc10))  xpc10 <= 13'sd501/*501:xpc10*/;
                  if ((13'sd502/*502:xpc10*/==xpc10))  xpc10 <= 13'sd503/*503:xpc10*/;
                  if ((13'sd503/*503:xpc10*/==xpc10))  xpc10 <= 13'sd504/*504:xpc10*/;
                  if ((13'sd504/*504:xpc10*/==xpc10))  xpc10 <= 13'sd505/*505:xpc10*/;
                  if ((13'sd506/*506:xpc10*/==xpc10))  xpc10 <= 13'sd507/*507:xpc10*/;
                  if ((13'sd507/*507:xpc10*/==xpc10))  xpc10 <= 13'sd508/*508:xpc10*/;
                  if ((13'sd508/*508:xpc10*/==xpc10))  xpc10 <= 13'sd509/*509:xpc10*/;
                  if ((13'sd510/*510:xpc10*/==xpc10))  xpc10 <= 13'sd511/*511:xpc10*/;
                  if ((13'sd511/*511:xpc10*/==xpc10))  xpc10 <= 13'sd512/*512:xpc10*/;
                  if ((13'sd512/*512:xpc10*/==xpc10))  xpc10 <= 13'sd513/*513:xpc10*/;
                  if ((13'sd516/*516:xpc10*/==xpc10))  xpc10 <= 13'sd517/*517:xpc10*/;
                  if ((13'sd517/*517:xpc10*/==xpc10))  xpc10 <= 13'sd518/*518:xpc10*/;
                  if ((13'sd518/*518:xpc10*/==xpc10))  xpc10 <= 13'sd519/*519:xpc10*/;
                  if ((13'sd519/*519:xpc10*/==xpc10))  xpc10 <= 13'sd520/*520:xpc10*/;
                  if ((13'sd521/*521:xpc10*/==xpc10))  xpc10 <= 13'sd522/*522:xpc10*/;
                  if ((13'sd527/*527:xpc10*/==xpc10))  xpc10 <= 13'sd528/*528:xpc10*/;
                  if ((13'sd528/*528:xpc10*/==xpc10))  xpc10 <= 13'sd529/*529:xpc10*/;
                  if ((13'sd529/*529:xpc10*/==xpc10))  xpc10 <= 13'sd530/*530:xpc10*/;
                  if ((13'sd531/*531:xpc10*/==xpc10))  xpc10 <= 13'sd532/*532:xpc10*/;
                  if ((13'sd532/*532:xpc10*/==xpc10))  xpc10 <= 13'sd533/*533:xpc10*/;
                  if ((13'sd533/*533:xpc10*/==xpc10))  xpc10 <= 13'sd534/*534:xpc10*/;
                  if ((13'sd538/*538:xpc10*/==xpc10))  xpc10 <= 13'sd539/*539:xpc10*/;
                  if ((13'sd539/*539:xpc10*/==xpc10))  xpc10 <= 13'sd540/*540:xpc10*/;
                  if ((13'sd540/*540:xpc10*/==xpc10))  xpc10 <= 13'sd541/*541:xpc10*/;
                  if ((13'sd542/*542:xpc10*/==xpc10))  xpc10 <= 13'sd543/*543:xpc10*/;
                  if ((13'sd543/*543:xpc10*/==xpc10))  xpc10 <= 13'sd544/*544:xpc10*/;
                  if ((13'sd544/*544:xpc10*/==xpc10))  xpc10 <= 13'sd545/*545:xpc10*/;
                  if ((13'sd548/*548:xpc10*/==xpc10))  xpc10 <= 13'sd549/*549:xpc10*/;
                  if ((13'sd549/*549:xpc10*/==xpc10))  xpc10 <= 13'sd550/*550:xpc10*/;
                  if ((13'sd550/*550:xpc10*/==xpc10))  xpc10 <= 13'sd551/*551:xpc10*/;
                  if ((13'sd552/*552:xpc10*/==xpc10))  xpc10 <= 13'sd553/*553:xpc10*/;
                  if ((13'sd553/*553:xpc10*/==xpc10))  xpc10 <= 13'sd554/*554:xpc10*/;
                  if ((13'sd554/*554:xpc10*/==xpc10))  xpc10 <= 13'sd555/*555:xpc10*/;
                  if ((13'sd556/*556:xpc10*/==xpc10))  xpc10 <= 13'sd557/*557:xpc10*/;
                  if ((13'sd557/*557:xpc10*/==xpc10))  xpc10 <= 13'sd558/*558:xpc10*/;
                  if ((13'sd558/*558:xpc10*/==xpc10))  xpc10 <= 13'sd559/*559:xpc10*/;
                  if ((13'sd560/*560:xpc10*/==xpc10))  xpc10 <= 13'sd561/*561:xpc10*/;
                  if ((13'sd561/*561:xpc10*/==xpc10))  xpc10 <= 13'sd562/*562:xpc10*/;
                  if ((13'sd562/*562:xpc10*/==xpc10))  xpc10 <= 13'sd563/*563:xpc10*/;
                  if ((13'sd566/*566:xpc10*/==xpc10))  xpc10 <= 13'sd567/*567:xpc10*/;
                  if ((13'sd567/*567:xpc10*/==xpc10))  xpc10 <= 13'sd568/*568:xpc10*/;
                  if ((13'sd568/*568:xpc10*/==xpc10))  xpc10 <= 13'sd569/*569:xpc10*/;
                  if ((13'sd570/*570:xpc10*/==xpc10))  xpc10 <= 13'sd571/*571:xpc10*/;
                  if ((13'sd571/*571:xpc10*/==xpc10))  xpc10 <= 13'sd572/*572:xpc10*/;
                  if ((13'sd572/*572:xpc10*/==xpc10))  xpc10 <= 13'sd573/*573:xpc10*/;
                  if ((13'sd576/*576:xpc10*/==xpc10))  xpc10 <= 13'sd577/*577:xpc10*/;
                  if ((13'sd577/*577:xpc10*/==xpc10))  xpc10 <= 13'sd578/*578:xpc10*/;
                  if ((13'sd578/*578:xpc10*/==xpc10))  xpc10 <= 13'sd579/*579:xpc10*/;
                  if ((13'sd580/*580:xpc10*/==xpc10))  xpc10 <= 13'sd581/*581:xpc10*/;
                  if ((13'sd581/*581:xpc10*/==xpc10))  xpc10 <= 13'sd582/*582:xpc10*/;
                  if ((13'sd582/*582:xpc10*/==xpc10))  xpc10 <= 13'sd583/*583:xpc10*/;
                  if ((13'sd587/*587:xpc10*/==xpc10))  xpc10 <= 13'sd588/*588:xpc10*/;
                  if ((13'sd588/*588:xpc10*/==xpc10))  xpc10 <= 13'sd589/*589:xpc10*/;
                  if ((13'sd589/*589:xpc10*/==xpc10))  xpc10 <= 13'sd590/*590:xpc10*/;
                  if ((13'sd590/*590:xpc10*/==xpc10))  xpc10 <= 13'sd591/*591:xpc10*/;
                  if ((13'sd591/*591:xpc10*/==xpc10))  xpc10 <= 13'sd592/*592:xpc10*/;
                  if ((13'sd592/*592:xpc10*/==xpc10))  xpc10 <= 13'sd593/*593:xpc10*/;
                  if ((13'sd593/*593:xpc10*/==xpc10))  xpc10 <= 13'sd594/*594:xpc10*/;
                  if ((13'sd595/*595:xpc10*/==xpc10))  xpc10 <= 13'sd596/*596:xpc10*/;
                  if ((13'sd596/*596:xpc10*/==xpc10))  xpc10 <= 13'sd597/*597:xpc10*/;
                  if ((13'sd597/*597:xpc10*/==xpc10))  xpc10 <= 13'sd598/*598:xpc10*/;
                  if ((13'sd599/*599:xpc10*/==xpc10))  xpc10 <= 13'sd600/*600:xpc10*/;
                  if ((13'sd600/*600:xpc10*/==xpc10))  xpc10 <= 13'sd601/*601:xpc10*/;
                  if ((13'sd601/*601:xpc10*/==xpc10))  xpc10 <= 13'sd602/*602:xpc10*/;
                  if ((13'sd603/*603:xpc10*/==xpc10))  xpc10 <= 13'sd604/*604:xpc10*/;
                  if ((13'sd604/*604:xpc10*/==xpc10))  xpc10 <= 13'sd605/*605:xpc10*/;
                  if ((13'sd605/*605:xpc10*/==xpc10))  xpc10 <= 13'sd606/*606:xpc10*/;
                  if ((13'sd607/*607:xpc10*/==xpc10))  xpc10 <= 13'sd608/*608:xpc10*/;
                  if ((13'sd608/*608:xpc10*/==xpc10))  xpc10 <= 13'sd609/*609:xpc10*/;
                  if ((13'sd609/*609:xpc10*/==xpc10))  xpc10 <= 13'sd610/*610:xpc10*/;
                  if ((13'sd611/*611:xpc10*/==xpc10))  xpc10 <= 13'sd612/*612:xpc10*/;
                  if ((13'sd612/*612:xpc10*/==xpc10))  xpc10 <= 13'sd613/*613:xpc10*/;
                  if ((13'sd613/*613:xpc10*/==xpc10))  xpc10 <= 13'sd614/*614:xpc10*/;
                  if ((13'sd615/*615:xpc10*/==xpc10))  xpc10 <= 13'sd616/*616:xpc10*/;
                  if ((13'sd621/*621:xpc10*/==xpc10))  xpc10 <= 13'sd622/*622:xpc10*/;
                  if ((13'sd622/*622:xpc10*/==xpc10))  xpc10 <= 13'sd623/*623:xpc10*/;
                  if ((13'sd623/*623:xpc10*/==xpc10))  xpc10 <= 13'sd624/*624:xpc10*/;
                  if ((13'sd625/*625:xpc10*/==xpc10))  xpc10 <= 13'sd626/*626:xpc10*/;
                  if ((13'sd626/*626:xpc10*/==xpc10))  xpc10 <= 13'sd627/*627:xpc10*/;
                  if ((13'sd627/*627:xpc10*/==xpc10))  xpc10 <= 13'sd628/*628:xpc10*/;
                  if ((13'sd632/*632:xpc10*/==xpc10))  xpc10 <= 13'sd633/*633:xpc10*/;
                  if ((13'sd633/*633:xpc10*/==xpc10))  xpc10 <= 13'sd634/*634:xpc10*/;
                  if ((13'sd634/*634:xpc10*/==xpc10))  xpc10 <= 13'sd635/*635:xpc10*/;
                  if ((13'sd636/*636:xpc10*/==xpc10))  xpc10 <= 13'sd637/*637:xpc10*/;
                  if ((13'sd637/*637:xpc10*/==xpc10))  xpc10 <= 13'sd638/*638:xpc10*/;
                  if ((13'sd638/*638:xpc10*/==xpc10))  xpc10 <= 13'sd639/*639:xpc10*/;
                  if ((13'sd642/*642:xpc10*/==xpc10))  xpc10 <= 13'sd643/*643:xpc10*/;
                  if ((13'sd643/*643:xpc10*/==xpc10))  xpc10 <= 13'sd644/*644:xpc10*/;
                  if ((13'sd644/*644:xpc10*/==xpc10))  xpc10 <= 13'sd645/*645:xpc10*/;
                  if ((13'sd646/*646:xpc10*/==xpc10))  xpc10 <= 13'sd647/*647:xpc10*/;
                  if ((13'sd647/*647:xpc10*/==xpc10))  xpc10 <= 13'sd648/*648:xpc10*/;
                  if ((13'sd648/*648:xpc10*/==xpc10))  xpc10 <= 13'sd649/*649:xpc10*/;
                  if ((13'sd650/*650:xpc10*/==xpc10))  xpc10 <= 13'sd651/*651:xpc10*/;
                  if ((13'sd651/*651:xpc10*/==xpc10))  xpc10 <= 13'sd652/*652:xpc10*/;
                  if ((13'sd652/*652:xpc10*/==xpc10))  xpc10 <= 13'sd653/*653:xpc10*/;
                  if ((13'sd654/*654:xpc10*/==xpc10))  xpc10 <= 13'sd655/*655:xpc10*/;
                  if ((13'sd655/*655:xpc10*/==xpc10))  xpc10 <= 13'sd656/*656:xpc10*/;
                  if ((13'sd656/*656:xpc10*/==xpc10))  xpc10 <= 13'sd657/*657:xpc10*/;
                  if ((13'sd660/*660:xpc10*/==xpc10))  xpc10 <= 13'sd661/*661:xpc10*/;
                  if ((13'sd661/*661:xpc10*/==xpc10))  xpc10 <= 13'sd662/*662:xpc10*/;
                  if ((13'sd662/*662:xpc10*/==xpc10))  xpc10 <= 13'sd663/*663:xpc10*/;
                  if ((13'sd664/*664:xpc10*/==xpc10))  xpc10 <= 13'sd665/*665:xpc10*/;
                  if ((13'sd665/*665:xpc10*/==xpc10))  xpc10 <= 13'sd666/*666:xpc10*/;
                  if ((13'sd666/*666:xpc10*/==xpc10))  xpc10 <= 13'sd667/*667:xpc10*/;
                  if ((13'sd670/*670:xpc10*/==xpc10))  xpc10 <= 13'sd671/*671:xpc10*/;
                  if ((13'sd671/*671:xpc10*/==xpc10))  xpc10 <= 13'sd672/*672:xpc10*/;
                  if ((13'sd672/*672:xpc10*/==xpc10))  xpc10 <= 13'sd673/*673:xpc10*/;
                  if ((13'sd674/*674:xpc10*/==xpc10))  xpc10 <= 13'sd675/*675:xpc10*/;
                  if ((13'sd675/*675:xpc10*/==xpc10))  xpc10 <= 13'sd676/*676:xpc10*/;
                  if ((13'sd676/*676:xpc10*/==xpc10))  xpc10 <= 13'sd677/*677:xpc10*/;
                  if ((13'sd681/*681:xpc10*/==xpc10))  xpc10 <= 13'sd682/*682:xpc10*/;
                  if ((13'sd682/*682:xpc10*/==xpc10))  xpc10 <= 13'sd683/*683:xpc10*/;
                  if ((13'sd683/*683:xpc10*/==xpc10))  xpc10 <= 13'sd684/*684:xpc10*/;
                  if ((13'sd684/*684:xpc10*/==xpc10))  xpc10 <= 13'sd685/*685:xpc10*/;
                  if ((13'sd685/*685:xpc10*/==xpc10))  xpc10 <= 13'sd686/*686:xpc10*/;
                  if ((13'sd686/*686:xpc10*/==xpc10))  xpc10 <= 13'sd687/*687:xpc10*/;
                  if ((13'sd687/*687:xpc10*/==xpc10))  xpc10 <= 13'sd688/*688:xpc10*/;
                  if ((13'sd689/*689:xpc10*/==xpc10))  xpc10 <= 13'sd690/*690:xpc10*/;
                  if ((13'sd690/*690:xpc10*/==xpc10))  xpc10 <= 13'sd691/*691:xpc10*/;
                  if ((13'sd691/*691:xpc10*/==xpc10))  xpc10 <= 13'sd692/*692:xpc10*/;
                  if ((13'sd693/*693:xpc10*/==xpc10))  xpc10 <= 13'sd694/*694:xpc10*/;
                  if ((13'sd694/*694:xpc10*/==xpc10))  xpc10 <= 13'sd695/*695:xpc10*/;
                  if ((13'sd695/*695:xpc10*/==xpc10))  xpc10 <= 13'sd696/*696:xpc10*/;
                  if ((13'sd697/*697:xpc10*/==xpc10))  xpc10 <= 13'sd698/*698:xpc10*/;
                  if ((13'sd698/*698:xpc10*/==xpc10))  xpc10 <= 13'sd699/*699:xpc10*/;
                  if ((13'sd699/*699:xpc10*/==xpc10))  xpc10 <= 13'sd700/*700:xpc10*/;
                  if ((13'sd701/*701:xpc10*/==xpc10))  xpc10 <= 13'sd702/*702:xpc10*/;
                  if ((13'sd702/*702:xpc10*/==xpc10))  xpc10 <= 13'sd703/*703:xpc10*/;
                  if ((13'sd703/*703:xpc10*/==xpc10))  xpc10 <= 13'sd704/*704:xpc10*/;
                  if ((13'sd705/*705:xpc10*/==xpc10))  xpc10 <= 13'sd706/*706:xpc10*/;
                  if ((13'sd706/*706:xpc10*/==xpc10))  xpc10 <= 13'sd707/*707:xpc10*/;
                  if ((13'sd707/*707:xpc10*/==xpc10))  xpc10 <= 13'sd708/*708:xpc10*/;
                  if ((13'sd711/*711:xpc10*/==xpc10))  xpc10 <= 13'sd712/*712:xpc10*/;
                  if ((13'sd712/*712:xpc10*/==xpc10))  xpc10 <= 13'sd713/*713:xpc10*/;
                  if ((13'sd713/*713:xpc10*/==xpc10))  xpc10 <= 13'sd714/*714:xpc10*/;
                  if ((13'sd715/*715:xpc10*/==xpc10))  xpc10 <= 13'sd716/*716:xpc10*/;
                  if ((13'sd716/*716:xpc10*/==xpc10))  xpc10 <= 13'sd717/*717:xpc10*/;
                  if ((13'sd717/*717:xpc10*/==xpc10))  xpc10 <= 13'sd718/*718:xpc10*/;
                  if ((13'sd722/*722:xpc10*/==xpc10))  xpc10 <= 13'sd723/*723:xpc10*/;
                  if ((13'sd723/*723:xpc10*/==xpc10))  xpc10 <= 13'sd724/*724:xpc10*/;
                  if ((13'sd724/*724:xpc10*/==xpc10))  xpc10 <= 13'sd725/*725:xpc10*/;
                  if ((13'sd726/*726:xpc10*/==xpc10))  xpc10 <= 13'sd727/*727:xpc10*/;
                  if ((13'sd727/*727:xpc10*/==xpc10))  xpc10 <= 13'sd728/*728:xpc10*/;
                  if ((13'sd728/*728:xpc10*/==xpc10))  xpc10 <= 13'sd729/*729:xpc10*/;
                  if ((13'sd732/*732:xpc10*/==xpc10))  xpc10 <= 13'sd733/*733:xpc10*/;
                  if ((13'sd733/*733:xpc10*/==xpc10))  xpc10 <= 13'sd734/*734:xpc10*/;
                  if ((13'sd734/*734:xpc10*/==xpc10))  xpc10 <= 13'sd735/*735:xpc10*/;
                  if ((13'sd736/*736:xpc10*/==xpc10))  xpc10 <= 13'sd737/*737:xpc10*/;
                  if ((13'sd737/*737:xpc10*/==xpc10))  xpc10 <= 13'sd738/*738:xpc10*/;
                  if ((13'sd738/*738:xpc10*/==xpc10))  xpc10 <= 13'sd739/*739:xpc10*/;
                  if ((13'sd742/*742:xpc10*/==xpc10))  xpc10 <= 13'sd743/*743:xpc10*/;
                  if ((13'sd743/*743:xpc10*/==xpc10))  xpc10 <= 13'sd744/*744:xpc10*/;
                  if ((13'sd744/*744:xpc10*/==xpc10))  xpc10 <= 13'sd745/*745:xpc10*/;
                  if ((13'sd746/*746:xpc10*/==xpc10))  xpc10 <= 13'sd747/*747:xpc10*/;
                  if ((13'sd747/*747:xpc10*/==xpc10))  xpc10 <= 13'sd748/*748:xpc10*/;
                  if ((13'sd748/*748:xpc10*/==xpc10))  xpc10 <= 13'sd749/*749:xpc10*/;
                  if ((13'sd752/*752:xpc10*/==xpc10))  xpc10 <= 13'sd753/*753:xpc10*/;
                  if ((13'sd753/*753:xpc10*/==xpc10))  xpc10 <= 13'sd754/*754:xpc10*/;
                  if ((13'sd754/*754:xpc10*/==xpc10))  xpc10 <= 13'sd755/*755:xpc10*/;
                  if ((13'sd756/*756:xpc10*/==xpc10))  xpc10 <= 13'sd757/*757:xpc10*/;
                  if ((13'sd757/*757:xpc10*/==xpc10))  xpc10 <= 13'sd758/*758:xpc10*/;
                  if ((13'sd758/*758:xpc10*/==xpc10))  xpc10 <= 13'sd759/*759:xpc10*/;
                  if ((13'sd763/*763:xpc10*/==xpc10))  xpc10 <= 13'sd764/*764:xpc10*/;
                  if ((13'sd764/*764:xpc10*/==xpc10))  xpc10 <= 13'sd765/*765:xpc10*/;
                  if ((13'sd765/*765:xpc10*/==xpc10))  xpc10 <= 13'sd766/*766:xpc10*/;
                  if ((13'sd766/*766:xpc10*/==xpc10))  xpc10 <= 13'sd767/*767:xpc10*/;
                  if ((13'sd767/*767:xpc10*/==xpc10))  xpc10 <= 13'sd768/*768:xpc10*/;
                  if ((13'sd768/*768:xpc10*/==xpc10))  xpc10 <= 13'sd769/*769:xpc10*/;
                  if ((13'sd769/*769:xpc10*/==xpc10))  xpc10 <= 13'sd770/*770:xpc10*/;
                  if ((13'sd771/*771:xpc10*/==xpc10))  xpc10 <= 13'sd772/*772:xpc10*/;
                  if ((13'sd772/*772:xpc10*/==xpc10))  xpc10 <= 13'sd773/*773:xpc10*/;
                  if ((13'sd773/*773:xpc10*/==xpc10))  xpc10 <= 13'sd774/*774:xpc10*/;
                  if ((13'sd775/*775:xpc10*/==xpc10))  xpc10 <= 13'sd776/*776:xpc10*/;
                  if ((13'sd776/*776:xpc10*/==xpc10))  xpc10 <= 13'sd777/*777:xpc10*/;
                  if ((13'sd777/*777:xpc10*/==xpc10))  xpc10 <= 13'sd778/*778:xpc10*/;
                  if ((13'sd779/*779:xpc10*/==xpc10))  xpc10 <= 13'sd780/*780:xpc10*/;
                  if ((13'sd780/*780:xpc10*/==xpc10))  xpc10 <= 13'sd781/*781:xpc10*/;
                  if ((13'sd781/*781:xpc10*/==xpc10))  xpc10 <= 13'sd782/*782:xpc10*/;
                  if ((13'sd784/*784:xpc10*/==xpc10))  xpc10 <= 13'sd785/*785:xpc10*/;
                  if ((13'sd785/*785:xpc10*/==xpc10))  xpc10 <= 13'sd786/*786:xpc10*/;
                  if ((13'sd786/*786:xpc10*/==xpc10))  xpc10 <= 13'sd787/*787:xpc10*/;
                  if ((13'sd788/*788:xpc10*/==xpc10))  xpc10 <= 13'sd789/*789:xpc10*/;
                  if ((13'sd789/*789:xpc10*/==xpc10))  xpc10 <= 13'sd790/*790:xpc10*/;
                  if ((13'sd790/*790:xpc10*/==xpc10))  xpc10 <= 13'sd791/*791:xpc10*/;
                  if ((13'sd793/*793:xpc10*/==xpc10))  xpc10 <= 13'sd794/*794:xpc10*/;
                  if ((13'sd794/*794:xpc10*/==xpc10))  xpc10 <= 13'sd795/*795:xpc10*/;
                  if ((13'sd795/*795:xpc10*/==xpc10))  xpc10 <= 13'sd796/*796:xpc10*/;
                  if ((13'sd797/*797:xpc10*/==xpc10))  xpc10 <= 13'sd798/*798:xpc10*/;
                  if ((13'sd798/*798:xpc10*/==xpc10))  xpc10 <= 13'sd799/*799:xpc10*/;
                  if ((13'sd799/*799:xpc10*/==xpc10))  xpc10 <= 13'sd800/*800:xpc10*/;
                  if ((13'sd802/*802:xpc10*/==xpc10))  xpc10 <= 13'sd803/*803:xpc10*/;
                  if ((13'sd803/*803:xpc10*/==xpc10))  xpc10 <= 13'sd804/*804:xpc10*/;
                  if ((13'sd804/*804:xpc10*/==xpc10))  xpc10 <= 13'sd805/*805:xpc10*/;
                  if ((13'sd813/*813:xpc10*/==xpc10))  xpc10 <= 13'sd814/*814:xpc10*/;
                  if ((13'sd814/*814:xpc10*/==xpc10))  xpc10 <= 13'sd815/*815:xpc10*/;
                  if ((13'sd815/*815:xpc10*/==xpc10))  xpc10 <= 13'sd816/*816:xpc10*/;
                  if ((13'sd817/*817:xpc10*/==xpc10))  xpc10 <= 13'sd818/*818:xpc10*/;
                  if ((13'sd818/*818:xpc10*/==xpc10))  xpc10 <= 13'sd819/*819:xpc10*/;
                  if ((13'sd819/*819:xpc10*/==xpc10))  xpc10 <= 13'sd820/*820:xpc10*/;
                  if ((13'sd821/*821:xpc10*/==xpc10))  xpc10 <= 13'sd822/*822:xpc10*/;
                  if ((13'sd822/*822:xpc10*/==xpc10))  xpc10 <= 13'sd823/*823:xpc10*/;
                  if ((13'sd823/*823:xpc10*/==xpc10))  xpc10 <= 13'sd824/*824:xpc10*/;
                  if ((13'sd827/*827:xpc10*/==xpc10))  xpc10 <= 13'sd828/*828:xpc10*/;
                  if ((13'sd828/*828:xpc10*/==xpc10))  xpc10 <= 13'sd829/*829:xpc10*/;
                  if ((13'sd829/*829:xpc10*/==xpc10))  xpc10 <= 13'sd830/*830:xpc10*/;
                  if ((13'sd831/*831:xpc10*/==xpc10))  xpc10 <= 13'sd832/*832:xpc10*/;
                  if ((13'sd832/*832:xpc10*/==xpc10))  xpc10 <= 13'sd833/*833:xpc10*/;
                  if ((13'sd833/*833:xpc10*/==xpc10))  xpc10 <= 13'sd834/*834:xpc10*/;
                  if ((13'sd837/*837:xpc10*/==xpc10))  xpc10 <= 13'sd838/*838:xpc10*/;
                  if ((13'sd838/*838:xpc10*/==xpc10))  xpc10 <= 13'sd839/*839:xpc10*/;
                  if ((13'sd839/*839:xpc10*/==xpc10))  xpc10 <= 13'sd840/*840:xpc10*/;
                  if ((13'sd841/*841:xpc10*/==xpc10))  xpc10 <= 13'sd842/*842:xpc10*/;
                  if ((13'sd842/*842:xpc10*/==xpc10))  xpc10 <= 13'sd843/*843:xpc10*/;
                  if ((13'sd843/*843:xpc10*/==xpc10))  xpc10 <= 13'sd844/*844:xpc10*/;
                  if ((13'sd848/*848:xpc10*/==xpc10))  xpc10 <= 13'sd849/*849:xpc10*/;
                  if ((13'sd849/*849:xpc10*/==xpc10))  xpc10 <= 13'sd850/*850:xpc10*/;
                  if ((13'sd850/*850:xpc10*/==xpc10))  xpc10 <= 13'sd851/*851:xpc10*/;
                  if ((13'sd851/*851:xpc10*/==xpc10))  xpc10 <= 13'sd852/*852:xpc10*/;
                  if ((13'sd852/*852:xpc10*/==xpc10))  xpc10 <= 13'sd853/*853:xpc10*/;
                  if ((13'sd853/*853:xpc10*/==xpc10))  xpc10 <= 13'sd854/*854:xpc10*/;
                  if ((13'sd854/*854:xpc10*/==xpc10))  xpc10 <= 13'sd855/*855:xpc10*/;
                  if ((13'sd856/*856:xpc10*/==xpc10))  xpc10 <= 13'sd857/*857:xpc10*/;
                  if ((13'sd857/*857:xpc10*/==xpc10))  xpc10 <= 13'sd858/*858:xpc10*/;
                  if ((13'sd858/*858:xpc10*/==xpc10))  xpc10 <= 13'sd859/*859:xpc10*/;
                  if ((13'sd860/*860:xpc10*/==xpc10))  xpc10 <= 13'sd861/*861:xpc10*/;
                  if ((13'sd861/*861:xpc10*/==xpc10))  xpc10 <= 13'sd862/*862:xpc10*/;
                  if ((13'sd862/*862:xpc10*/==xpc10))  xpc10 <= 13'sd863/*863:xpc10*/;
                  if ((13'sd864/*864:xpc10*/==xpc10))  xpc10 <= 13'sd865/*865:xpc10*/;
                  if ((13'sd865/*865:xpc10*/==xpc10))  xpc10 <= 13'sd866/*866:xpc10*/;
                  if ((13'sd866/*866:xpc10*/==xpc10))  xpc10 <= 13'sd867/*867:xpc10*/;
                  if ((13'sd868/*868:xpc10*/==xpc10))  xpc10 <= 13'sd869/*869:xpc10*/;
                  if ((13'sd869/*869:xpc10*/==xpc10))  xpc10 <= 13'sd870/*870:xpc10*/;
                  if ((13'sd870/*870:xpc10*/==xpc10))  xpc10 <= 13'sd871/*871:xpc10*/;
                  if ((13'sd873/*873:xpc10*/==xpc10))  xpc10 <= 13'sd874/*874:xpc10*/;
                  if ((13'sd875/*875:xpc10*/==xpc10))  xpc10 <= 13'sd876/*876:xpc10*/;
                  if ((13'sd876/*876:xpc10*/==xpc10))  xpc10 <= 13'sd877/*877:xpc10*/;
                  if ((13'sd877/*877:xpc10*/==xpc10))  xpc10 <= 13'sd878/*878:xpc10*/;
                  if ((13'sd879/*879:xpc10*/==xpc10))  xpc10 <= 13'sd880/*880:xpc10*/;
                  if ((13'sd880/*880:xpc10*/==xpc10))  xpc10 <= 13'sd881/*881:xpc10*/;
                  if ((13'sd881/*881:xpc10*/==xpc10))  xpc10 <= 13'sd882/*882:xpc10*/;
                  if ((13'sd883/*883:xpc10*/==xpc10))  xpc10 <= 13'sd884/*884:xpc10*/;
                  if ((13'sd884/*884:xpc10*/==xpc10))  xpc10 <= 13'sd885/*885:xpc10*/;
                  if ((13'sd885/*885:xpc10*/==xpc10))  xpc10 <= 13'sd886/*886:xpc10*/;
                  if ((13'sd886/*886:xpc10*/==xpc10))  xpc10 <= 13'sd887/*887:xpc10*/;
                  if ((13'sd888/*888:xpc10*/==xpc10))  xpc10 <= 13'sd889/*889:xpc10*/;
                  if ((13'sd889/*889:xpc10*/==xpc10))  xpc10 <= 13'sd890/*890:xpc10*/;
                  if ((13'sd890/*890:xpc10*/==xpc10))  xpc10 <= 13'sd891/*891:xpc10*/;
                  if ((13'sd892/*892:xpc10*/==xpc10))  xpc10 <= 13'sd893/*893:xpc10*/;
                  if ((13'sd893/*893:xpc10*/==xpc10))  xpc10 <= 13'sd894/*894:xpc10*/;
                  if ((13'sd894/*894:xpc10*/==xpc10))  xpc10 <= 13'sd895/*895:xpc10*/;
                  if ((13'sd896/*896:xpc10*/==xpc10))  xpc10 <= 13'sd897/*897:xpc10*/;
                  if ((13'sd897/*897:xpc10*/==xpc10))  xpc10 <= 13'sd898/*898:xpc10*/;
                  if ((13'sd902/*902:xpc10*/==xpc10))  xpc10 <= 13'sd903/*903:xpc10*/;
                  if ((13'sd903/*903:xpc10*/==xpc10))  xpc10 <= 13'sd904/*904:xpc10*/;
                  if ((13'sd904/*904:xpc10*/==xpc10))  xpc10 <= 13'sd905/*905:xpc10*/;
                  if ((13'sd907/*907:xpc10*/==xpc10))  xpc10 <= 13'sd908/*908:xpc10*/;
                  if ((13'sd908/*908:xpc10*/==xpc10))  xpc10 <= 13'sd909/*909:xpc10*/;
                  if ((13'sd909/*909:xpc10*/==xpc10))  xpc10 <= 13'sd910/*910:xpc10*/;
                  if ((13'sd911/*911:xpc10*/==xpc10))  xpc10 <= 13'sd912/*912:xpc10*/;
                  if ((13'sd913/*913:xpc10*/==xpc10))  xpc10 <= 13'sd914/*914:xpc10*/;
                  if ((13'sd915/*915:xpc10*/==xpc10))  xpc10 <= 13'sd916/*916:xpc10*/;
                  if ((13'sd916/*916:xpc10*/==xpc10))  xpc10 <= 13'sd917/*917:xpc10*/;
                  if ((13'sd917/*917:xpc10*/==xpc10))  xpc10 <= 13'sd918/*918:xpc10*/;
                  if ((13'sd919/*919:xpc10*/==xpc10))  xpc10 <= 13'sd920/*920:xpc10*/;
                  if ((13'sd920/*920:xpc10*/==xpc10))  xpc10 <= 13'sd921/*921:xpc10*/;
                  if ((13'sd921/*921:xpc10*/==xpc10))  xpc10 <= 13'sd922/*922:xpc10*/;
                  if ((13'sd922/*922:xpc10*/==xpc10))  xpc10 <= 13'sd923/*923:xpc10*/;
                  if ((13'sd924/*924:xpc10*/==xpc10))  xpc10 <= 13'sd925/*925:xpc10*/;
                  if ((13'sd925/*925:xpc10*/==xpc10))  xpc10 <= 13'sd926/*926:xpc10*/;
                  if ((13'sd926/*926:xpc10*/==xpc10))  xpc10 <= 13'sd927/*927:xpc10*/;
                  if ((13'sd928/*928:xpc10*/==xpc10))  xpc10 <= 13'sd929/*929:xpc10*/;
                  if ((13'sd929/*929:xpc10*/==xpc10))  xpc10 <= 13'sd930/*930:xpc10*/;
                  if ((13'sd930/*930:xpc10*/==xpc10))  xpc10 <= 13'sd931/*931:xpc10*/;
                  if ((13'sd931/*931:xpc10*/==xpc10))  xpc10 <= 13'sd932/*932:xpc10*/;
                  if ((13'sd933/*933:xpc10*/==xpc10))  xpc10 <= 13'sd934/*934:xpc10*/;
                  if ((13'sd935/*935:xpc10*/==xpc10))  xpc10 <= 13'sd936/*936:xpc10*/;
                  if ((13'sd936/*936:xpc10*/==xpc10))  xpc10 <= 13'sd937/*937:xpc10*/;
                  if ((13'sd937/*937:xpc10*/==xpc10))  xpc10 <= 13'sd938/*938:xpc10*/;
                  if ((13'sd939/*939:xpc10*/==xpc10))  xpc10 <= 13'sd940/*940:xpc10*/;
                  if ((13'sd940/*940:xpc10*/==xpc10))  xpc10 <= 13'sd941/*941:xpc10*/;
                  if ((13'sd941/*941:xpc10*/==xpc10))  xpc10 <= 13'sd942/*942:xpc10*/;
                  if ((13'sd942/*942:xpc10*/==xpc10))  xpc10 <= 13'sd943/*943:xpc10*/;
                  if ((13'sd944/*944:xpc10*/==xpc10))  xpc10 <= 13'sd945/*945:xpc10*/;
                  if ((13'sd946/*946:xpc10*/==xpc10))  xpc10 <= 13'sd947/*947:xpc10*/;
                  if ((13'sd947/*947:xpc10*/==xpc10))  xpc10 <= 13'sd948/*948:xpc10*/;
                  if ((13'sd949/*949:xpc10*/==xpc10))  xpc10 <= 13'sd950/*950:xpc10*/;
                  if ((13'sd950/*950:xpc10*/==xpc10))  xpc10 <= 13'sd951/*951:xpc10*/;
                  if ((13'sd952/*952:xpc10*/==xpc10))  xpc10 <= 13'sd953/*953:xpc10*/;
                  if ((13'sd953/*953:xpc10*/==xpc10))  xpc10 <= 13'sd941/*941:xpc10*/;
                  if ((13'sd954/*954:xpc10*/==xpc10))  xpc10 <= 13'sd955/*955:xpc10*/;
                  if ((13'sd955/*955:xpc10*/==xpc10))  xpc10 <= 13'sd956/*956:xpc10*/;
                  if ((13'sd958/*958:xpc10*/==xpc10))  xpc10 <= 13'sd908/*908:xpc10*/;
                  if ((13'sd959/*959:xpc10*/==xpc10))  xpc10 <= 13'sd960/*960:xpc10*/;
                  if ((13'sd960/*960:xpc10*/==xpc10))  xpc10 <= 13'sd961/*961:xpc10*/;
                  if ((13'sd961/*961:xpc10*/==xpc10))  xpc10 <= 13'sd962/*962:xpc10*/;
                  if ((13'sd962/*962:xpc10*/==xpc10))  xpc10 <= 13'sd963/*963:xpc10*/;
                  if ((13'sd963/*963:xpc10*/==xpc10))  xpc10 <= 13'sd964/*964:xpc10*/;
                  if ((13'sd965/*965:xpc10*/==xpc10))  xpc10 <= 13'sd966/*966:xpc10*/;
                  if ((13'sd966/*966:xpc10*/==xpc10))  xpc10 <= 13'sd967/*967:xpc10*/;
                  if ((13'sd967/*967:xpc10*/==xpc10))  xpc10 <= 13'sd968/*968:xpc10*/;
                  if ((13'sd970/*970:xpc10*/==xpc10))  xpc10 <= 13'sd971/*971:xpc10*/;
                  if ((13'sd971/*971:xpc10*/==xpc10))  xpc10 <= 13'sd972/*972:xpc10*/;
                  if ((13'sd972/*972:xpc10*/==xpc10))  xpc10 <= 13'sd973/*973:xpc10*/;
                  if ((13'sd974/*974:xpc10*/==xpc10))  xpc10 <= 13'sd975/*975:xpc10*/;
                  if ((13'sd975/*975:xpc10*/==xpc10))  xpc10 <= 13'sd976/*976:xpc10*/;
                  if ((13'sd976/*976:xpc10*/==xpc10))  xpc10 <= 13'sd977/*977:xpc10*/;
                  if ((13'sd979/*979:xpc10*/==xpc10))  xpc10 <= 13'sd980/*980:xpc10*/;
                  if ((13'sd980/*980:xpc10*/==xpc10))  xpc10 <= 13'sd981/*981:xpc10*/;
                  if ((13'sd981/*981:xpc10*/==xpc10))  xpc10 <= 13'sd982/*982:xpc10*/;
                  if ((13'sd983/*983:xpc10*/==xpc10))  xpc10 <= 13'sd984/*984:xpc10*/;
                  if ((13'sd984/*984:xpc10*/==xpc10))  xpc10 <= 13'sd985/*985:xpc10*/;
                  if ((13'sd985/*985:xpc10*/==xpc10))  xpc10 <= 13'sd986/*986:xpc10*/;
                  if ((13'sd987/*987:xpc10*/==xpc10))  xpc10 <= 13'sd988/*988:xpc10*/;
                  if ((13'sd988/*988:xpc10*/==xpc10))  xpc10 <= 13'sd989/*989:xpc10*/;
                  if ((13'sd989/*989:xpc10*/==xpc10))  xpc10 <= 13'sd990/*990:xpc10*/;
                  if ((13'sd991/*991:xpc10*/==xpc10))  xpc10 <= 13'sd889/*889:xpc10*/;
                  if ((13'sd992/*992:xpc10*/==xpc10))  xpc10 <= 13'sd993/*993:xpc10*/;
                  if ((13'sd993/*993:xpc10*/==xpc10))  xpc10 <= 13'sd994/*994:xpc10*/;
                  if ((13'sd995/*995:xpc10*/==xpc10))  xpc10 <= 13'sd988/*988:xpc10*/;
                  if ((13'sd996/*996:xpc10*/==xpc10))  xpc10 <= 13'sd997/*997:xpc10*/;
                  if ((13'sd997/*997:xpc10*/==xpc10))  xpc10 <= 13'sd998/*998:xpc10*/;
                  if ((13'sd999/*999:xpc10*/==xpc10))  xpc10 <= 13'sd1000/*1000:xpc10*/;
                  if ((13'sd1000/*1000:xpc10*/==xpc10))  xpc10 <= 13'sd1001/*1001:xpc10*/;
                  if ((13'sd1001/*1001:xpc10*/==xpc10))  xpc10 <= 13'sd1002/*1002:xpc10*/;
                  if ((13'sd1003/*1003:xpc10*/==xpc10))  xpc10 <= 13'sd1004/*1004:xpc10*/;
                  if ((13'sd1004/*1004:xpc10*/==xpc10))  xpc10 <= 13'sd1005/*1005:xpc10*/;
                  if ((13'sd1005/*1005:xpc10*/==xpc10))  xpc10 <= 13'sd1006/*1006:xpc10*/;
                  if ((13'sd1007/*1007:xpc10*/==xpc10))  xpc10 <= 13'sd889/*889:xpc10*/;
                  if ((13'sd1008/*1008:xpc10*/==xpc10))  xpc10 <= 13'sd1009/*1009:xpc10*/;
                  if ((13'sd1009/*1009:xpc10*/==xpc10))  xpc10 <= 13'sd1010/*1010:xpc10*/;
                  if ((13'sd1011/*1011:xpc10*/==xpc10))  xpc10 <= 13'sd1004/*1004:xpc10*/;
                  if ((13'sd1012/*1012:xpc10*/==xpc10))  xpc10 <= 13'sd1013/*1013:xpc10*/;
                  if ((13'sd1013/*1013:xpc10*/==xpc10))  xpc10 <= 13'sd1014/*1014:xpc10*/;
                  if ((13'sd1015/*1015:xpc10*/==xpc10))  xpc10 <= 13'sd975/*975:xpc10*/;
                  if ((13'sd1016/*1016:xpc10*/==xpc10))  xpc10 <= 13'sd1017/*1017:xpc10*/;
                  if ((13'sd1017/*1017:xpc10*/==xpc10))  xpc10 <= 13'sd1018/*1018:xpc10*/;
                  if ((13'sd1019/*1019:xpc10*/==xpc10))  xpc10 <= 13'sd1020/*1020:xpc10*/;
                  if ((13'sd1020/*1020:xpc10*/==xpc10))  xpc10 <= 13'sd1021/*1021:xpc10*/;
                  if ((13'sd1021/*1021:xpc10*/==xpc10))  xpc10 <= 13'sd1022/*1022:xpc10*/;
                  if ((13'sd1023/*1023:xpc10*/==xpc10))  xpc10 <= 13'sd861/*861:xpc10*/;
                  if ((13'sd1024/*1024:xpc10*/==xpc10))  xpc10 <= 13'sd1025/*1025:xpc10*/;
                  if ((13'sd1025/*1025:xpc10*/==xpc10))  xpc10 <= 13'sd1026/*1026:xpc10*/;
                  if ((13'sd1027/*1027:xpc10*/==xpc10))  xpc10 <= 13'sd1028/*1028:xpc10*/;
                  if ((13'sd1028/*1028:xpc10*/==xpc10))  xpc10 <= 13'sd1029/*1029:xpc10*/;
                  if ((13'sd1029/*1029:xpc10*/==xpc10))  xpc10 <= 13'sd1030/*1030:xpc10*/;
                  if ((13'sd1031/*1031:xpc10*/==xpc10))  xpc10 <= 13'sd861/*861:xpc10*/;
                  if ((13'sd1032/*1032:xpc10*/==xpc10))  xpc10 <= 13'sd1033/*1033:xpc10*/;
                  if ((13'sd1033/*1033:xpc10*/==xpc10))  xpc10 <= 13'sd1034/*1034:xpc10*/;
                  if ((13'sd1035/*1035:xpc10*/==xpc10))  xpc10 <= 13'sd861/*861:xpc10*/;
                  if ((13'sd1036/*1036:xpc10*/==xpc10))  xpc10 <= 13'sd1037/*1037:xpc10*/;
                  if ((13'sd1037/*1037:xpc10*/==xpc10))  xpc10 <= 13'sd1038/*1038:xpc10*/;
                  if ((13'sd1039/*1039:xpc10*/==xpc10))  xpc10 <= 13'sd842/*842:xpc10*/;
                  if ((13'sd1040/*1040:xpc10*/==xpc10))  xpc10 <= 13'sd1041/*1041:xpc10*/;
                  if ((13'sd1041/*1041:xpc10*/==xpc10))  xpc10 <= 13'sd1042/*1042:xpc10*/;
                  if ((13'sd1043/*1043:xpc10*/==xpc10))  xpc10 <= 13'sd832/*832:xpc10*/;
                  if ((13'sd1044/*1044:xpc10*/==xpc10))  xpc10 <= 13'sd1045/*1045:xpc10*/;
                  if ((13'sd1045/*1045:xpc10*/==xpc10))  xpc10 <= 13'sd1046/*1046:xpc10*/;
                  if ((13'sd1047/*1047:xpc10*/==xpc10))  xpc10 <= 13'sd865/*865:xpc10*/;
                  if ((13'sd1048/*1048:xpc10*/==xpc10))  xpc10 <= 13'sd1049/*1049:xpc10*/;
                  if ((13'sd1049/*1049:xpc10*/==xpc10))  xpc10 <= 13'sd1050/*1050:xpc10*/;
                  if ((13'sd1051/*1051:xpc10*/==xpc10))  xpc10 <= 13'sd1052/*1052:xpc10*/;
                  if ((13'sd1052/*1052:xpc10*/==xpc10))  xpc10 <= 13'sd1053/*1053:xpc10*/;
                  if ((13'sd1053/*1053:xpc10*/==xpc10))  xpc10 <= 13'sd1054/*1054:xpc10*/;
                  if ((13'sd1055/*1055:xpc10*/==xpc10))  xpc10 <= 13'sd1056/*1056:xpc10*/;
                  if ((13'sd1056/*1056:xpc10*/==xpc10))  xpc10 <= 13'sd1057/*1057:xpc10*/;
                  if ((13'sd1057/*1057:xpc10*/==xpc10))  xpc10 <= 13'sd1058/*1058:xpc10*/;
                  if ((13'sd1059/*1059:xpc10*/==xpc10))  xpc10 <= 13'sd1060/*1060:xpc10*/;
                  if ((13'sd1060/*1060:xpc10*/==xpc10))  xpc10 <= 13'sd1061/*1061:xpc10*/;
                  if ((13'sd1061/*1061:xpc10*/==xpc10))  xpc10 <= 13'sd1062/*1062:xpc10*/;
                  if ((13'sd1063/*1063:xpc10*/==xpc10))  xpc10 <= 13'sd1064/*1064:xpc10*/;
                  if ((13'sd1064/*1064:xpc10*/==xpc10))  xpc10 <= 13'sd1065/*1065:xpc10*/;
                  if ((13'sd1065/*1065:xpc10*/==xpc10))  xpc10 <= 13'sd1066/*1066:xpc10*/;
                  if ((13'sd1068/*1068:xpc10*/==xpc10))  xpc10 <= 13'sd1069/*1069:xpc10*/;
                  if ((13'sd1069/*1069:xpc10*/==xpc10))  xpc10 <= 13'sd1070/*1070:xpc10*/;
                  if ((13'sd1070/*1070:xpc10*/==xpc10))  xpc10 <= 13'sd1071/*1071:xpc10*/;
                  if ((13'sd1075/*1075:xpc10*/==xpc10))  xpc10 <= 13'sd1076/*1076:xpc10*/;
                  if ((13'sd1076/*1076:xpc10*/==xpc10))  xpc10 <= 13'sd1077/*1077:xpc10*/;
                  if ((13'sd1077/*1077:xpc10*/==xpc10))  xpc10 <= 13'sd1078/*1078:xpc10*/;
                  if ((13'sd1080/*1080:xpc10*/==xpc10))  xpc10 <= 13'sd1081/*1081:xpc10*/;
                  if ((13'sd1081/*1081:xpc10*/==xpc10))  xpc10 <= 13'sd1082/*1082:xpc10*/;
                  if ((13'sd1082/*1082:xpc10*/==xpc10))  xpc10 <= 13'sd1083/*1083:xpc10*/;
                  if ((13'sd1085/*1085:xpc10*/==xpc10))  xpc10 <= 13'sd1086/*1086:xpc10*/;
                  if ((13'sd1086/*1086:xpc10*/==xpc10))  xpc10 <= 13'sd1087/*1087:xpc10*/;
                  if ((13'sd1088/*1088:xpc10*/==xpc10))  xpc10 <= 13'sd1089/*1089:xpc10*/;
                  if ((13'sd1089/*1089:xpc10*/==xpc10))  xpc10 <= 13'sd1090/*1090:xpc10*/;
                  if ((13'sd1090/*1090:xpc10*/==xpc10))  xpc10 <= 13'sd1091/*1091:xpc10*/;
                  if ((13'sd1093/*1093:xpc10*/==xpc10))  xpc10 <= 13'sd1094/*1094:xpc10*/;
                  if ((13'sd1094/*1094:xpc10*/==xpc10))  xpc10 <= 13'sd1095/*1095:xpc10*/;
                  if ((13'sd1095/*1095:xpc10*/==xpc10))  xpc10 <= 13'sd1096/*1096:xpc10*/;
                  if ((13'sd1097/*1097:xpc10*/==xpc10))  xpc10 <= 13'sd1098/*1098:xpc10*/;
                  if ((13'sd1098/*1098:xpc10*/==xpc10))  xpc10 <= 13'sd1099/*1099:xpc10*/;
                  if ((13'sd1099/*1099:xpc10*/==xpc10))  xpc10 <= 13'sd1100/*1100:xpc10*/;
                  if ((13'sd1101/*1101:xpc10*/==xpc10))  xpc10 <= 13'sd1102/*1102:xpc10*/;
                  if ((13'sd1102/*1102:xpc10*/==xpc10))  xpc10 <= 13'sd1103/*1103:xpc10*/;
                  if ((13'sd1103/*1103:xpc10*/==xpc10))  xpc10 <= 13'sd1104/*1104:xpc10*/;
                  if ((13'sd1105/*1105:xpc10*/==xpc10))  xpc10 <= 13'sd1106/*1106:xpc10*/;
                  if ((13'sd1106/*1106:xpc10*/==xpc10))  xpc10 <= 13'sd1107/*1107:xpc10*/;
                  if ((13'sd1107/*1107:xpc10*/==xpc10))  xpc10 <= 13'sd1108/*1108:xpc10*/;
                  if ((13'sd1108/*1108:xpc10*/==xpc10))  xpc10 <= 13'sd1109/*1109:xpc10*/;
                  if ((13'sd1110/*1110:xpc10*/==xpc10))  xpc10 <= 13'sd1111/*1111:xpc10*/;
                  if ((13'sd1111/*1111:xpc10*/==xpc10))  xpc10 <= 13'sd1112/*1112:xpc10*/;
                  if ((13'sd1112/*1112:xpc10*/==xpc10))  xpc10 <= 13'sd1113/*1113:xpc10*/;
                  if ((13'sd1114/*1114:xpc10*/==xpc10))  xpc10 <= 13'sd1115/*1115:xpc10*/;
                  if ((13'sd1115/*1115:xpc10*/==xpc10))  xpc10 <= 13'sd1116/*1116:xpc10*/;
                  if ((13'sd1116/*1116:xpc10*/==xpc10))  xpc10 <= 13'sd1117/*1117:xpc10*/;
                  if ((13'sd1121/*1121:xpc10*/==xpc10))  xpc10 <= 13'sd1122/*1122:xpc10*/;
                  if ((13'sd1122/*1122:xpc10*/==xpc10))  xpc10 <= 13'sd1123/*1123:xpc10*/;
                  if ((13'sd1123/*1123:xpc10*/==xpc10))  xpc10 <= 13'sd1124/*1124:xpc10*/;
                  if ((13'sd1126/*1126:xpc10*/==xpc10))  xpc10 <= 13'sd1127/*1127:xpc10*/;
                  if ((13'sd1127/*1127:xpc10*/==xpc10))  xpc10 <= 13'sd1128/*1128:xpc10*/;
                  if ((13'sd1128/*1128:xpc10*/==xpc10))  xpc10 <= 13'sd1129/*1129:xpc10*/;
                  if ((13'sd1130/*1130:xpc10*/==xpc10))  xpc10 <= 13'sd1131/*1131:xpc10*/;
                  if ((13'sd1131/*1131:xpc10*/==xpc10))  xpc10 <= 13'sd1132/*1132:xpc10*/;
                  if ((13'sd1132/*1132:xpc10*/==xpc10))  xpc10 <= 13'sd1133/*1133:xpc10*/;
                  if ((13'sd1134/*1134:xpc10*/==xpc10))  xpc10 <= 13'sd865/*865:xpc10*/;
                  if ((13'sd1135/*1135:xpc10*/==xpc10))  xpc10 <= 13'sd1136/*1136:xpc10*/;
                  if ((13'sd1136/*1136:xpc10*/==xpc10))  xpc10 <= 13'sd1137/*1137:xpc10*/;
                  if ((13'sd1139/*1139:xpc10*/==xpc10))  xpc10 <= 13'sd1127/*1127:xpc10*/;
                  if ((13'sd1140/*1140:xpc10*/==xpc10))  xpc10 <= 13'sd1141/*1141:xpc10*/;
                  if ((13'sd1141/*1141:xpc10*/==xpc10))  xpc10 <= 13'sd1142/*1142:xpc10*/;
                  if ((13'sd1143/*1143:xpc10*/==xpc10))  xpc10 <= 13'sd1115/*1115:xpc10*/;
                  if ((13'sd1144/*1144:xpc10*/==xpc10))  xpc10 <= 13'sd1145/*1145:xpc10*/;
                  if ((13'sd1145/*1145:xpc10*/==xpc10))  xpc10 <= 13'sd1146/*1146:xpc10*/;
                  if ((13'sd1147/*1147:xpc10*/==xpc10))  xpc10 <= 13'sd1148/*1148:xpc10*/;
                  if ((13'sd1148/*1148:xpc10*/==xpc10))  xpc10 <= 13'sd1149/*1149:xpc10*/;
                  if ((13'sd1149/*1149:xpc10*/==xpc10))  xpc10 <= 13'sd1150/*1150:xpc10*/;
                  if ((13'sd1150/*1150:xpc10*/==xpc10))  xpc10 <= 13'sd1151/*1151:xpc10*/;
                  if ((13'sd1152/*1152:xpc10*/==xpc10))  xpc10 <= 13'sd1153/*1153:xpc10*/;
                  if ((13'sd1153/*1153:xpc10*/==xpc10))  xpc10 <= 13'sd1154/*1154:xpc10*/;
                  if ((13'sd1154/*1154:xpc10*/==xpc10))  xpc10 <= 13'sd1155/*1155:xpc10*/;
                  if ((13'sd1156/*1156:xpc10*/==xpc10))  xpc10 <= 13'sd1157/*1157:xpc10*/;
                  if ((13'sd1157/*1157:xpc10*/==xpc10))  xpc10 <= 13'sd1158/*1158:xpc10*/;
                  if ((13'sd1158/*1158:xpc10*/==xpc10))  xpc10 <= 13'sd1159/*1159:xpc10*/;
                  if ((13'sd1162/*1162:xpc10*/==xpc10))  xpc10 <= 13'sd1163/*1163:xpc10*/;
                  if ((13'sd1163/*1163:xpc10*/==xpc10))  xpc10 <= 13'sd1164/*1164:xpc10*/;
                  if ((13'sd1164/*1164:xpc10*/==xpc10))  xpc10 <= 13'sd1165/*1165:xpc10*/;
                  if ((13'sd1166/*1166:xpc10*/==xpc10))  xpc10 <= 13'sd1167/*1167:xpc10*/;
                  if ((13'sd1167/*1167:xpc10*/==xpc10))  xpc10 <= 13'sd1168/*1168:xpc10*/;
                  if ((13'sd1168/*1168:xpc10*/==xpc10))  xpc10 <= 13'sd1169/*1169:xpc10*/;
                  if ((13'sd1169/*1169:xpc10*/==xpc10))  xpc10 <= 13'sd1170/*1170:xpc10*/;
                  if ((13'sd1170/*1170:xpc10*/==xpc10))  xpc10 <= 13'sd1171/*1171:xpc10*/;
                  if ((13'sd1171/*1171:xpc10*/==xpc10))  xpc10 <= 13'sd1172/*1172:xpc10*/;
                  if ((13'sd1172/*1172:xpc10*/==xpc10))  xpc10 <= 13'sd1173/*1173:xpc10*/;
                  if ((13'sd1174/*1174:xpc10*/==xpc10))  xpc10 <= 13'sd1175/*1175:xpc10*/;
                  if ((13'sd1175/*1175:xpc10*/==xpc10))  xpc10 <= 13'sd1176/*1176:xpc10*/;
                  if ((13'sd1176/*1176:xpc10*/==xpc10))  xpc10 <= 13'sd1177/*1177:xpc10*/;
                  if ((13'sd1177/*1177:xpc10*/==xpc10))  xpc10 <= 13'sd1178/*1178:xpc10*/;
                  if ((13'sd1178/*1178:xpc10*/==xpc10))  xpc10 <= 13'sd1179/*1179:xpc10*/;
                  if ((13'sd1179/*1179:xpc10*/==xpc10))  xpc10 <= 13'sd1180/*1180:xpc10*/;
                  if ((13'sd1180/*1180:xpc10*/==xpc10))  xpc10 <= 13'sd1181/*1181:xpc10*/;
                  if ((13'sd1183/*1183:xpc10*/==xpc10))  xpc10 <= 13'sd1184/*1184:xpc10*/;
                  if ((13'sd1184/*1184:xpc10*/==xpc10))  xpc10 <= 13'sd1185/*1185:xpc10*/;
                  if ((13'sd1185/*1185:xpc10*/==xpc10))  xpc10 <= 13'sd1186/*1186:xpc10*/;
                  if ((13'sd1187/*1187:xpc10*/==xpc10))  xpc10 <= 13'sd1188/*1188:xpc10*/;
                  if ((13'sd1188/*1188:xpc10*/==xpc10))  xpc10 <= 13'sd1189/*1189:xpc10*/;
                  if ((13'sd1189/*1189:xpc10*/==xpc10))  xpc10 <= 13'sd1190/*1190:xpc10*/;
                  if ((13'sd1191/*1191:xpc10*/==xpc10))  xpc10 <= 13'sd1192/*1192:xpc10*/;
                  if ((13'sd1192/*1192:xpc10*/==xpc10))  xpc10 <= 13'sd1193/*1193:xpc10*/;
                  if ((13'sd1193/*1193:xpc10*/==xpc10))  xpc10 <= 13'sd1194/*1194:xpc10*/;
                  if ((13'sd1195/*1195:xpc10*/==xpc10))  xpc10 <= 13'sd1196/*1196:xpc10*/;
                  if ((13'sd1196/*1196:xpc10*/==xpc10))  xpc10 <= 13'sd1197/*1197:xpc10*/;
                  if ((13'sd1197/*1197:xpc10*/==xpc10))  xpc10 <= 13'sd1198/*1198:xpc10*/;
                  if ((13'sd1199/*1199:xpc10*/==xpc10))  xpc10 <= 13'sd1200/*1200:xpc10*/;
                  if ((13'sd1200/*1200:xpc10*/==xpc10))  xpc10 <= 13'sd1201/*1201:xpc10*/;
                  if ((13'sd1201/*1201:xpc10*/==xpc10))  xpc10 <= 13'sd1202/*1202:xpc10*/;
                  if ((13'sd1203/*1203:xpc10*/==xpc10))  xpc10 <= 13'sd1204/*1204:xpc10*/;
                  if ((13'sd1204/*1204:xpc10*/==xpc10))  xpc10 <= 13'sd1205/*1205:xpc10*/;
                  if ((13'sd1205/*1205:xpc10*/==xpc10))  xpc10 <= 13'sd1206/*1206:xpc10*/;
                  if ((13'sd1207/*1207:xpc10*/==xpc10))  xpc10 <= 13'sd1131/*1131:xpc10*/;
                  if ((13'sd1208/*1208:xpc10*/==xpc10))  xpc10 <= 13'sd1209/*1209:xpc10*/;
                  if ((13'sd1209/*1209:xpc10*/==xpc10))  xpc10 <= 13'sd1210/*1210:xpc10*/;
                  if ((13'sd1211/*1211:xpc10*/==xpc10))  xpc10 <= 13'sd1204/*1204:xpc10*/;
                  if ((13'sd1212/*1212:xpc10*/==xpc10))  xpc10 <= 13'sd1213/*1213:xpc10*/;
                  if ((13'sd1213/*1213:xpc10*/==xpc10))  xpc10 <= 13'sd1214/*1214:xpc10*/;
                  if ((13'sd1215/*1215:xpc10*/==xpc10))  xpc10 <= 13'sd1216/*1216:xpc10*/;
                  if ((13'sd1216/*1216:xpc10*/==xpc10))  xpc10 <= 13'sd1217/*1217:xpc10*/;
                  if ((13'sd1217/*1217:xpc10*/==xpc10))  xpc10 <= 13'sd1218/*1218:xpc10*/;
                  if ((13'sd1222/*1222:xpc10*/==xpc10))  xpc10 <= 13'sd1223/*1223:xpc10*/;
                  if ((13'sd1223/*1223:xpc10*/==xpc10))  xpc10 <= 13'sd1224/*1224:xpc10*/;
                  if ((13'sd1224/*1224:xpc10*/==xpc10))  xpc10 <= 13'sd1225/*1225:xpc10*/;
                  if ((13'sd1227/*1227:xpc10*/==xpc10))  xpc10 <= 13'sd1228/*1228:xpc10*/;
                  if ((13'sd1228/*1228:xpc10*/==xpc10))  xpc10 <= 13'sd1229/*1229:xpc10*/;
                  if ((13'sd1229/*1229:xpc10*/==xpc10))  xpc10 <= 13'sd1230/*1230:xpc10*/;
                  if ((13'sd1231/*1231:xpc10*/==xpc10))  xpc10 <= 13'sd1157/*1157:xpc10*/;
                  if ((13'sd1232/*1232:xpc10*/==xpc10))  xpc10 <= 13'sd1233/*1233:xpc10*/;
                  if ((13'sd1233/*1233:xpc10*/==xpc10))  xpc10 <= 13'sd1234/*1234:xpc10*/;
                  if ((13'sd1236/*1236:xpc10*/==xpc10))  xpc10 <= 13'sd1228/*1228:xpc10*/;
                  if ((13'sd1237/*1237:xpc10*/==xpc10))  xpc10 <= 13'sd1238/*1238:xpc10*/;
                  if ((13'sd1238/*1238:xpc10*/==xpc10))  xpc10 <= 13'sd1239/*1239:xpc10*/;
                  if ((13'sd1240/*1240:xpc10*/==xpc10))  xpc10 <= 13'sd1241/*1241:xpc10*/;
                  if ((13'sd1241/*1241:xpc10*/==xpc10))  xpc10 <= 13'sd1242/*1242:xpc10*/;
                  if ((13'sd1242/*1242:xpc10*/==xpc10))  xpc10 <= 13'sd1243/*1243:xpc10*/;
                  if ((13'sd1244/*1244:xpc10*/==xpc10))  xpc10 <= 13'sd1245/*1245:xpc10*/;
                  if ((13'sd1245/*1245:xpc10*/==xpc10))  xpc10 <= 13'sd1246/*1246:xpc10*/;
                  if ((13'sd1246/*1246:xpc10*/==xpc10))  xpc10 <= 13'sd1247/*1247:xpc10*/;
                  if ((13'sd1248/*1248:xpc10*/==xpc10))  xpc10 <= 13'sd1157/*1157:xpc10*/;
                  if ((13'sd1249/*1249:xpc10*/==xpc10))  xpc10 <= 13'sd1250/*1250:xpc10*/;
                  if ((13'sd1250/*1250:xpc10*/==xpc10))  xpc10 <= 13'sd1251/*1251:xpc10*/;
                  if ((13'sd1252/*1252:xpc10*/==xpc10))  xpc10 <= 13'sd1245/*1245:xpc10*/;
                  if ((13'sd1253/*1253:xpc10*/==xpc10))  xpc10 <= 13'sd1254/*1254:xpc10*/;
                  if ((13'sd1254/*1254:xpc10*/==xpc10))  xpc10 <= 13'sd1255/*1255:xpc10*/;
                  if ((13'sd1256/*1256:xpc10*/==xpc10))  xpc10 <= 13'sd1257/*1257:xpc10*/;
                  if ((13'sd1257/*1257:xpc10*/==xpc10))  xpc10 <= 13'sd1258/*1258:xpc10*/;
                  if ((13'sd1258/*1258:xpc10*/==xpc10))  xpc10 <= 13'sd1259/*1259:xpc10*/;
                  if ((13'sd1263/*1263:xpc10*/==xpc10))  xpc10 <= 13'sd1264/*1264:xpc10*/;
                  if ((13'sd1264/*1264:xpc10*/==xpc10))  xpc10 <= 13'sd1265/*1265:xpc10*/;
                  if ((13'sd1265/*1265:xpc10*/==xpc10))  xpc10 <= 13'sd1266/*1266:xpc10*/;
                  if ((13'sd1268/*1268:xpc10*/==xpc10))  xpc10 <= 13'sd1269/*1269:xpc10*/;
                  if ((13'sd1269/*1269:xpc10*/==xpc10))  xpc10 <= 13'sd1270/*1270:xpc10*/;
                  if ((13'sd1270/*1270:xpc10*/==xpc10))  xpc10 <= 13'sd1271/*1271:xpc10*/;
                  if ((13'sd1272/*1272:xpc10*/==xpc10))  xpc10 <= 13'sd1064/*1064:xpc10*/;
                  if ((13'sd1273/*1273:xpc10*/==xpc10))  xpc10 <= 13'sd1274/*1274:xpc10*/;
                  if ((13'sd1274/*1274:xpc10*/==xpc10))  xpc10 <= 13'sd1275/*1275:xpc10*/;
                  if ((13'sd1277/*1277:xpc10*/==xpc10))  xpc10 <= 13'sd1269/*1269:xpc10*/;
                  if ((13'sd1278/*1278:xpc10*/==xpc10))  xpc10 <= 13'sd1279/*1279:xpc10*/;
                  if ((13'sd1279/*1279:xpc10*/==xpc10))  xpc10 <= 13'sd1280/*1280:xpc10*/;
                  if ((13'sd1281/*1281:xpc10*/==xpc10))  xpc10 <= 13'sd1282/*1282:xpc10*/;
                  if ((13'sd1282/*1282:xpc10*/==xpc10))  xpc10 <= 13'sd1283/*1283:xpc10*/;
                  if ((13'sd1283/*1283:xpc10*/==xpc10))  xpc10 <= 13'sd1284/*1284:xpc10*/;
                  if ((13'sd1285/*1285:xpc10*/==xpc10))  xpc10 <= 13'sd1286/*1286:xpc10*/;
                  if ((13'sd1286/*1286:xpc10*/==xpc10))  xpc10 <= 13'sd1287/*1287:xpc10*/;
                  if ((13'sd1287/*1287:xpc10*/==xpc10))  xpc10 <= 13'sd1288/*1288:xpc10*/;
                  if ((13'sd1289/*1289:xpc10*/==xpc10))  xpc10 <= 13'sd1064/*1064:xpc10*/;
                  if ((13'sd1290/*1290:xpc10*/==xpc10))  xpc10 <= 13'sd1291/*1291:xpc10*/;
                  if ((13'sd1291/*1291:xpc10*/==xpc10))  xpc10 <= 13'sd1292/*1292:xpc10*/;
                  if ((13'sd1293/*1293:xpc10*/==xpc10))  xpc10 <= 13'sd1286/*1286:xpc10*/;
                  if ((13'sd1294/*1294:xpc10*/==xpc10))  xpc10 <= 13'sd1295/*1295:xpc10*/;
                  if ((13'sd1295/*1295:xpc10*/==xpc10))  xpc10 <= 13'sd1296/*1296:xpc10*/;
                  if ((13'sd1297/*1297:xpc10*/==xpc10))  xpc10 <= 13'sd1056/*1056:xpc10*/;
                  if ((13'sd1298/*1298:xpc10*/==xpc10))  xpc10 <= 13'sd1299/*1299:xpc10*/;
                  if ((13'sd1299/*1299:xpc10*/==xpc10))  xpc10 <= 13'sd1300/*1300:xpc10*/;
                  if ((13'sd1301/*1301:xpc10*/==xpc10))  xpc10 <= 13'sd1302/*1302:xpc10*/;
                  if ((13'sd1302/*1302:xpc10*/==xpc10))  xpc10 <= 13'sd1303/*1303:xpc10*/;
                  if ((13'sd1303/*1303:xpc10*/==xpc10))  xpc10 <= 13'sd1304/*1304:xpc10*/;
                  if ((13'sd1305/*1305:xpc10*/==xpc10))  xpc10 <= 13'sd1306/*1306:xpc10*/;
                  if ((13'sd1306/*1306:xpc10*/==xpc10))  xpc10 <= 13'sd1307/*1307:xpc10*/;
                  if ((13'sd1307/*1307:xpc10*/==xpc10))  xpc10 <= 13'sd1308/*1308:xpc10*/;
                  if ((13'sd1309/*1309:xpc10*/==xpc10))  xpc10 <= 13'sd1310/*1310:xpc10*/;
                  if ((13'sd1310/*1310:xpc10*/==xpc10))  xpc10 <= 13'sd1311/*1311:xpc10*/;
                  if ((13'sd1311/*1311:xpc10*/==xpc10))  xpc10 <= 13'sd1312/*1312:xpc10*/;
                  if ((13'sd1315/*1315:xpc10*/==xpc10))  xpc10 <= 13'sd1316/*1316:xpc10*/;
                  if ((13'sd1316/*1316:xpc10*/==xpc10))  xpc10 <= 13'sd1317/*1317:xpc10*/;
                  if ((13'sd1317/*1317:xpc10*/==xpc10))  xpc10 <= 13'sd1318/*1318:xpc10*/;
                  if ((13'sd1319/*1319:xpc10*/==xpc10))  xpc10 <= 13'sd1320/*1320:xpc10*/;
                  if ((13'sd1320/*1320:xpc10*/==xpc10))  xpc10 <= 13'sd1321/*1321:xpc10*/;
                  if ((13'sd1321/*1321:xpc10*/==xpc10))  xpc10 <= 13'sd1322/*1322:xpc10*/;
                  if ((13'sd1325/*1325:xpc10*/==xpc10))  xpc10 <= 13'sd1326/*1326:xpc10*/;
                  if ((13'sd1326/*1326:xpc10*/==xpc10))  xpc10 <= 13'sd1327/*1327:xpc10*/;
                  if ((13'sd1327/*1327:xpc10*/==xpc10))  xpc10 <= 13'sd1328/*1328:xpc10*/;
                  if ((13'sd1329/*1329:xpc10*/==xpc10))  xpc10 <= 13'sd1330/*1330:xpc10*/;
                  if ((13'sd1330/*1330:xpc10*/==xpc10))  xpc10 <= 13'sd1331/*1331:xpc10*/;
                  if ((13'sd1331/*1331:xpc10*/==xpc10))  xpc10 <= 13'sd1332/*1332:xpc10*/;
                  if ((13'sd1336/*1336:xpc10*/==xpc10))  xpc10 <= 13'sd1337/*1337:xpc10*/;
                  if ((13'sd1337/*1337:xpc10*/==xpc10))  xpc10 <= 13'sd1338/*1338:xpc10*/;
                  if ((13'sd1338/*1338:xpc10*/==xpc10))  xpc10 <= 13'sd1339/*1339:xpc10*/;
                  if ((13'sd1339/*1339:xpc10*/==xpc10))  xpc10 <= 13'sd1340/*1340:xpc10*/;
                  if ((13'sd1340/*1340:xpc10*/==xpc10))  xpc10 <= 13'sd1341/*1341:xpc10*/;
                  if ((13'sd1341/*1341:xpc10*/==xpc10))  xpc10 <= 13'sd1342/*1342:xpc10*/;
                  if ((13'sd1342/*1342:xpc10*/==xpc10))  xpc10 <= 13'sd1343/*1343:xpc10*/;
                  if ((13'sd1344/*1344:xpc10*/==xpc10))  xpc10 <= 13'sd1345/*1345:xpc10*/;
                  if ((13'sd1345/*1345:xpc10*/==xpc10))  xpc10 <= 13'sd1346/*1346:xpc10*/;
                  if ((13'sd1346/*1346:xpc10*/==xpc10))  xpc10 <= 13'sd1347/*1347:xpc10*/;
                  if ((13'sd1348/*1348:xpc10*/==xpc10))  xpc10 <= 13'sd1349/*1349:xpc10*/;
                  if ((13'sd1349/*1349:xpc10*/==xpc10))  xpc10 <= 13'sd1350/*1350:xpc10*/;
                  if ((13'sd1350/*1350:xpc10*/==xpc10))  xpc10 <= 13'sd1351/*1351:xpc10*/;
                  if ((13'sd1352/*1352:xpc10*/==xpc10))  xpc10 <= 13'sd865/*865:xpc10*/;
                  if ((13'sd1353/*1353:xpc10*/==xpc10))  xpc10 <= 13'sd1354/*1354:xpc10*/;
                  if ((13'sd1354/*1354:xpc10*/==xpc10))  xpc10 <= 13'sd1355/*1355:xpc10*/;
                  if ((13'sd1356/*1356:xpc10*/==xpc10))  xpc10 <= 13'sd1357/*1357:xpc10*/;
                  if ((13'sd1357/*1357:xpc10*/==xpc10))  xpc10 <= 13'sd1358/*1358:xpc10*/;
                  if ((13'sd1358/*1358:xpc10*/==xpc10))  xpc10 <= 13'sd1359/*1359:xpc10*/;
                  if ((13'sd1360/*1360:xpc10*/==xpc10))  xpc10 <= 13'sd1349/*1349:xpc10*/;
                  if ((13'sd1361/*1361:xpc10*/==xpc10))  xpc10 <= 13'sd1362/*1362:xpc10*/;
                  if ((13'sd1362/*1362:xpc10*/==xpc10))  xpc10 <= 13'sd1363/*1363:xpc10*/;
                  if ((13'sd1364/*1364:xpc10*/==xpc10))  xpc10 <= 13'sd1365/*1365:xpc10*/;
                  if ((13'sd1365/*1365:xpc10*/==xpc10))  xpc10 <= 13'sd1366/*1366:xpc10*/;
                  if ((13'sd1366/*1366:xpc10*/==xpc10))  xpc10 <= 13'sd1367/*1367:xpc10*/;
                  if ((13'sd1368/*1368:xpc10*/==xpc10))  xpc10 <= 13'sd1349/*1349:xpc10*/;
                  if ((13'sd1369/*1369:xpc10*/==xpc10))  xpc10 <= 13'sd1370/*1370:xpc10*/;
                  if ((13'sd1370/*1370:xpc10*/==xpc10))  xpc10 <= 13'sd1371/*1371:xpc10*/;
                  if ((13'sd1372/*1372:xpc10*/==xpc10))  xpc10 <= 13'sd1349/*1349:xpc10*/;
                  if ((13'sd1373/*1373:xpc10*/==xpc10))  xpc10 <= 13'sd1374/*1374:xpc10*/;
                  if ((13'sd1374/*1374:xpc10*/==xpc10))  xpc10 <= 13'sd1375/*1375:xpc10*/;
                  if ((13'sd1376/*1376:xpc10*/==xpc10))  xpc10 <= 13'sd1330/*1330:xpc10*/;
                  if ((13'sd1377/*1377:xpc10*/==xpc10))  xpc10 <= 13'sd1378/*1378:xpc10*/;
                  if ((13'sd1378/*1378:xpc10*/==xpc10))  xpc10 <= 13'sd1379/*1379:xpc10*/;
                  if ((13'sd1380/*1380:xpc10*/==xpc10))  xpc10 <= 13'sd1320/*1320:xpc10*/;
                  if ((13'sd1381/*1381:xpc10*/==xpc10))  xpc10 <= 13'sd1382/*1382:xpc10*/;
                  if ((13'sd1382/*1382:xpc10*/==xpc10))  xpc10 <= 13'sd1383/*1383:xpc10*/;
                  if ((13'sd1384/*1384:xpc10*/==xpc10))  xpc10 <= 13'sd1385/*1385:xpc10*/;
                  if ((13'sd1385/*1385:xpc10*/==xpc10))  xpc10 <= 13'sd1386/*1386:xpc10*/;
                  if ((13'sd1386/*1386:xpc10*/==xpc10))  xpc10 <= 13'sd1387/*1387:xpc10*/;
                  if ((13'sd1388/*1388:xpc10*/==xpc10))  xpc10 <= 13'sd1389/*1389:xpc10*/;
                  if ((13'sd1389/*1389:xpc10*/==xpc10))  xpc10 <= 13'sd1390/*1390:xpc10*/;
                  if ((13'sd1390/*1390:xpc10*/==xpc10))  xpc10 <= 13'sd1391/*1391:xpc10*/;
                  if ((13'sd1392/*1392:xpc10*/==xpc10))  xpc10 <= 13'sd865/*865:xpc10*/;
                  if ((13'sd1393/*1393:xpc10*/==xpc10))  xpc10 <= 13'sd1394/*1394:xpc10*/;
                  if ((13'sd1394/*1394:xpc10*/==xpc10))  xpc10 <= 13'sd1395/*1395:xpc10*/;
                  if ((13'sd1396/*1396:xpc10*/==xpc10))  xpc10 <= 13'sd1389/*1389:xpc10*/;
                  if ((13'sd1397/*1397:xpc10*/==xpc10))  xpc10 <= 13'sd1398/*1398:xpc10*/;
                  if ((13'sd1398/*1398:xpc10*/==xpc10))  xpc10 <= 13'sd1399/*1399:xpc10*/;
                  if ((13'sd1400/*1400:xpc10*/==xpc10))  xpc10 <= 13'sd1401/*1401:xpc10*/;
                  if ((13'sd1401/*1401:xpc10*/==xpc10))  xpc10 <= 13'sd1402/*1402:xpc10*/;
                  if ((13'sd1402/*1402:xpc10*/==xpc10))  xpc10 <= 13'sd1403/*1403:xpc10*/;
                  if ((13'sd1404/*1404:xpc10*/==xpc10))  xpc10 <= 13'sd1405/*1405:xpc10*/;
                  if ((13'sd1405/*1405:xpc10*/==xpc10))  xpc10 <= 13'sd1406/*1406:xpc10*/;
                  if ((13'sd1406/*1406:xpc10*/==xpc10))  xpc10 <= 13'sd1407/*1407:xpc10*/;
                  if ((13'sd1408/*1408:xpc10*/==xpc10))  xpc10 <= 13'sd1409/*1409:xpc10*/;
                  if ((13'sd1409/*1409:xpc10*/==xpc10))  xpc10 <= 13'sd1410/*1410:xpc10*/;
                  if ((13'sd1410/*1410:xpc10*/==xpc10))  xpc10 <= 13'sd1411/*1411:xpc10*/;
                  if ((13'sd1412/*1412:xpc10*/==xpc10))  xpc10 <= 13'sd1413/*1413:xpc10*/;
                  if ((13'sd1413/*1413:xpc10*/==xpc10))  xpc10 <= 13'sd1414/*1414:xpc10*/;
                  if ((13'sd1414/*1414:xpc10*/==xpc10))  xpc10 <= 13'sd1415/*1415:xpc10*/;
                  if ((13'sd1417/*1417:xpc10*/==xpc10))  xpc10 <= 13'sd1069/*1069:xpc10*/;
                  if ((13'sd1418/*1418:xpc10*/==xpc10))  xpc10 <= 13'sd1419/*1419:xpc10*/;
                  if ((13'sd1419/*1419:xpc10*/==xpc10))  xpc10 <= 13'sd1420/*1420:xpc10*/;
                  if ((13'sd1421/*1421:xpc10*/==xpc10))  xpc10 <= 13'sd1422/*1422:xpc10*/;
                  if ((13'sd1422/*1422:xpc10*/==xpc10))  xpc10 <= 13'sd1423/*1423:xpc10*/;
                  if ((13'sd1423/*1423:xpc10*/==xpc10))  xpc10 <= 13'sd1424/*1424:xpc10*/;
                  if ((13'sd1428/*1428:xpc10*/==xpc10))  xpc10 <= 13'sd1429/*1429:xpc10*/;
                  if ((13'sd1429/*1429:xpc10*/==xpc10))  xpc10 <= 13'sd1430/*1430:xpc10*/;
                  if ((13'sd1430/*1430:xpc10*/==xpc10))  xpc10 <= 13'sd1431/*1431:xpc10*/;
                  if ((13'sd1433/*1433:xpc10*/==xpc10))  xpc10 <= 13'sd1434/*1434:xpc10*/;
                  if ((13'sd1434/*1434:xpc10*/==xpc10))  xpc10 <= 13'sd1435/*1435:xpc10*/;
                  if ((13'sd1435/*1435:xpc10*/==xpc10))  xpc10 <= 13'sd1436/*1436:xpc10*/;
                  if ((13'sd1437/*1437:xpc10*/==xpc10))  xpc10 <= 13'sd1413/*1413:xpc10*/;
                  if ((13'sd1438/*1438:xpc10*/==xpc10))  xpc10 <= 13'sd1439/*1439:xpc10*/;
                  if ((13'sd1439/*1439:xpc10*/==xpc10))  xpc10 <= 13'sd1440/*1440:xpc10*/;
                  if ((13'sd1442/*1442:xpc10*/==xpc10))  xpc10 <= 13'sd1434/*1434:xpc10*/;
                  if ((13'sd1443/*1443:xpc10*/==xpc10))  xpc10 <= 13'sd1444/*1444:xpc10*/;
                  if ((13'sd1444/*1444:xpc10*/==xpc10))  xpc10 <= 13'sd1445/*1445:xpc10*/;
                  if ((13'sd1446/*1446:xpc10*/==xpc10))  xpc10 <= 13'sd1447/*1447:xpc10*/;
                  if ((13'sd1447/*1447:xpc10*/==xpc10))  xpc10 <= 13'sd1448/*1448:xpc10*/;
                  if ((13'sd1448/*1448:xpc10*/==xpc10))  xpc10 <= 13'sd1449/*1449:xpc10*/;
                  if ((13'sd1450/*1450:xpc10*/==xpc10))  xpc10 <= 13'sd1451/*1451:xpc10*/;
                  if ((13'sd1451/*1451:xpc10*/==xpc10))  xpc10 <= 13'sd1452/*1452:xpc10*/;
                  if ((13'sd1452/*1452:xpc10*/==xpc10))  xpc10 <= 13'sd1453/*1453:xpc10*/;
                  if ((13'sd1454/*1454:xpc10*/==xpc10))  xpc10 <= 13'sd1413/*1413:xpc10*/;
                  if ((13'sd1455/*1455:xpc10*/==xpc10))  xpc10 <= 13'sd1456/*1456:xpc10*/;
                  if ((13'sd1456/*1456:xpc10*/==xpc10))  xpc10 <= 13'sd1457/*1457:xpc10*/;
                  if ((13'sd1458/*1458:xpc10*/==xpc10))  xpc10 <= 13'sd1451/*1451:xpc10*/;
                  if ((13'sd1459/*1459:xpc10*/==xpc10))  xpc10 <= 13'sd1460/*1460:xpc10*/;
                  if ((13'sd1460/*1460:xpc10*/==xpc10))  xpc10 <= 13'sd1461/*1461:xpc10*/;
                  if ((13'sd1462/*1462:xpc10*/==xpc10))  xpc10 <= 13'sd1405/*1405:xpc10*/;
                  if ((13'sd1463/*1463:xpc10*/==xpc10))  xpc10 <= 13'sd1464/*1464:xpc10*/;
                  if ((13'sd1464/*1464:xpc10*/==xpc10))  xpc10 <= 13'sd1465/*1465:xpc10*/;
                  if ((13'sd1466/*1466:xpc10*/==xpc10))  xpc10 <= 13'sd1467/*1467:xpc10*/;
                  if ((13'sd1467/*1467:xpc10*/==xpc10))  xpc10 <= 13'sd1468/*1468:xpc10*/;
                  if ((13'sd1468/*1468:xpc10*/==xpc10))  xpc10 <= 13'sd1469/*1469:xpc10*/;
                  if ((13'sd1470/*1470:xpc10*/==xpc10))  xpc10 <= 13'sd1471/*1471:xpc10*/;
                  if ((13'sd1471/*1471:xpc10*/==xpc10))  xpc10 <= 13'sd1472/*1472:xpc10*/;
                  if ((13'sd1472/*1472:xpc10*/==xpc10))  xpc10 <= 13'sd1473/*1473:xpc10*/;
                  if ((13'sd1474/*1474:xpc10*/==xpc10))  xpc10 <= 13'sd1475/*1475:xpc10*/;
                  if ((13'sd1475/*1475:xpc10*/==xpc10))  xpc10 <= 13'sd1476/*1476:xpc10*/;
                  if ((13'sd1476/*1476:xpc10*/==xpc10))  xpc10 <= 13'sd1477/*1477:xpc10*/;
                  if ((13'sd1480/*1480:xpc10*/==xpc10))  xpc10 <= 13'sd1481/*1481:xpc10*/;
                  if ((13'sd1481/*1481:xpc10*/==xpc10))  xpc10 <= 13'sd1482/*1482:xpc10*/;
                  if ((13'sd1482/*1482:xpc10*/==xpc10))  xpc10 <= 13'sd1483/*1483:xpc10*/;
                  if ((13'sd1484/*1484:xpc10*/==xpc10))  xpc10 <= 13'sd1485/*1485:xpc10*/;
                  if ((13'sd1485/*1485:xpc10*/==xpc10))  xpc10 <= 13'sd1486/*1486:xpc10*/;
                  if ((13'sd1486/*1486:xpc10*/==xpc10))  xpc10 <= 13'sd1487/*1487:xpc10*/;
                  if ((13'sd1490/*1490:xpc10*/==xpc10))  xpc10 <= 13'sd1491/*1491:xpc10*/;
                  if ((13'sd1491/*1491:xpc10*/==xpc10))  xpc10 <= 13'sd1492/*1492:xpc10*/;
                  if ((13'sd1492/*1492:xpc10*/==xpc10))  xpc10 <= 13'sd1493/*1493:xpc10*/;
                  if ((13'sd1494/*1494:xpc10*/==xpc10))  xpc10 <= 13'sd1495/*1495:xpc10*/;
                  if ((13'sd1495/*1495:xpc10*/==xpc10))  xpc10 <= 13'sd1496/*1496:xpc10*/;
                  if ((13'sd1496/*1496:xpc10*/==xpc10))  xpc10 <= 13'sd1497/*1497:xpc10*/;
                  if ((13'sd1501/*1501:xpc10*/==xpc10))  xpc10 <= 13'sd1502/*1502:xpc10*/;
                  if ((13'sd1502/*1502:xpc10*/==xpc10))  xpc10 <= 13'sd1503/*1503:xpc10*/;
                  if ((13'sd1503/*1503:xpc10*/==xpc10))  xpc10 <= 13'sd1504/*1504:xpc10*/;
                  if ((13'sd1504/*1504:xpc10*/==xpc10))  xpc10 <= 13'sd1505/*1505:xpc10*/;
                  if ((13'sd1505/*1505:xpc10*/==xpc10))  xpc10 <= 13'sd1506/*1506:xpc10*/;
                  if ((13'sd1506/*1506:xpc10*/==xpc10))  xpc10 <= 13'sd1507/*1507:xpc10*/;
                  if ((13'sd1507/*1507:xpc10*/==xpc10))  xpc10 <= 13'sd1508/*1508:xpc10*/;
                  if ((13'sd1509/*1509:xpc10*/==xpc10))  xpc10 <= 13'sd1510/*1510:xpc10*/;
                  if ((13'sd1510/*1510:xpc10*/==xpc10))  xpc10 <= 13'sd1511/*1511:xpc10*/;
                  if ((13'sd1511/*1511:xpc10*/==xpc10))  xpc10 <= 13'sd1512/*1512:xpc10*/;
                  if ((13'sd1513/*1513:xpc10*/==xpc10))  xpc10 <= 13'sd1514/*1514:xpc10*/;
                  if ((13'sd1514/*1514:xpc10*/==xpc10))  xpc10 <= 13'sd1515/*1515:xpc10*/;
                  if ((13'sd1515/*1515:xpc10*/==xpc10))  xpc10 <= 13'sd1516/*1516:xpc10*/;
                  if ((13'sd1517/*1517:xpc10*/==xpc10))  xpc10 <= 13'sd865/*865:xpc10*/;
                  if ((13'sd1518/*1518:xpc10*/==xpc10))  xpc10 <= 13'sd1519/*1519:xpc10*/;
                  if ((13'sd1519/*1519:xpc10*/==xpc10))  xpc10 <= 13'sd1520/*1520:xpc10*/;
                  if ((13'sd1521/*1521:xpc10*/==xpc10))  xpc10 <= 13'sd1522/*1522:xpc10*/;
                  if ((13'sd1522/*1522:xpc10*/==xpc10))  xpc10 <= 13'sd1523/*1523:xpc10*/;
                  if ((13'sd1523/*1523:xpc10*/==xpc10))  xpc10 <= 13'sd1524/*1524:xpc10*/;
                  if ((13'sd1525/*1525:xpc10*/==xpc10))  xpc10 <= 13'sd1514/*1514:xpc10*/;
                  if ((13'sd1526/*1526:xpc10*/==xpc10))  xpc10 <= 13'sd1527/*1527:xpc10*/;
                  if ((13'sd1527/*1527:xpc10*/==xpc10))  xpc10 <= 13'sd1528/*1528:xpc10*/;
                  if ((13'sd1529/*1529:xpc10*/==xpc10))  xpc10 <= 13'sd1530/*1530:xpc10*/;
                  if ((13'sd1530/*1530:xpc10*/==xpc10))  xpc10 <= 13'sd1531/*1531:xpc10*/;
                  if ((13'sd1531/*1531:xpc10*/==xpc10))  xpc10 <= 13'sd1532/*1532:xpc10*/;
                  if ((13'sd1533/*1533:xpc10*/==xpc10))  xpc10 <= 13'sd1514/*1514:xpc10*/;
                  if ((13'sd1534/*1534:xpc10*/==xpc10))  xpc10 <= 13'sd1535/*1535:xpc10*/;
                  if ((13'sd1535/*1535:xpc10*/==xpc10))  xpc10 <= 13'sd1536/*1536:xpc10*/;
                  if ((13'sd1537/*1537:xpc10*/==xpc10))  xpc10 <= 13'sd1514/*1514:xpc10*/;
                  if ((13'sd1538/*1538:xpc10*/==xpc10))  xpc10 <= 13'sd1539/*1539:xpc10*/;
                  if ((13'sd1539/*1539:xpc10*/==xpc10))  xpc10 <= 13'sd1540/*1540:xpc10*/;
                  if ((13'sd1541/*1541:xpc10*/==xpc10))  xpc10 <= 13'sd1495/*1495:xpc10*/;
                  if ((13'sd1542/*1542:xpc10*/==xpc10))  xpc10 <= 13'sd1543/*1543:xpc10*/;
                  if ((13'sd1543/*1543:xpc10*/==xpc10))  xpc10 <= 13'sd1544/*1544:xpc10*/;
                  if ((13'sd1545/*1545:xpc10*/==xpc10))  xpc10 <= 13'sd1485/*1485:xpc10*/;
                  if ((13'sd1546/*1546:xpc10*/==xpc10))  xpc10 <= 13'sd1547/*1547:xpc10*/;
                  if ((13'sd1547/*1547:xpc10*/==xpc10))  xpc10 <= 13'sd1548/*1548:xpc10*/;
                  if ((13'sd1549/*1549:xpc10*/==xpc10))  xpc10 <= 13'sd865/*865:xpc10*/;
                  if ((13'sd1550/*1550:xpc10*/==xpc10))  xpc10 <= 13'sd1551/*1551:xpc10*/;
                  if ((13'sd1551/*1551:xpc10*/==xpc10))  xpc10 <= 13'sd1552/*1552:xpc10*/;
                  if ((13'sd1553/*1553:xpc10*/==xpc10))  xpc10 <= 13'sd1554/*1554:xpc10*/;
                  if ((13'sd1554/*1554:xpc10*/==xpc10))  xpc10 <= 13'sd1555/*1555:xpc10*/;
                  if ((13'sd1555/*1555:xpc10*/==xpc10))  xpc10 <= 13'sd1556/*1556:xpc10*/;
                  if ((13'sd1557/*1557:xpc10*/==xpc10))  xpc10 <= 13'sd1558/*1558:xpc10*/;
                  if ((13'sd1558/*1558:xpc10*/==xpc10))  xpc10 <= 13'sd1559/*1559:xpc10*/;
                  if ((13'sd1559/*1559:xpc10*/==xpc10))  xpc10 <= 13'sd1560/*1560:xpc10*/;
                  if ((13'sd1561/*1561:xpc10*/==xpc10))  xpc10 <= 13'sd1562/*1562:xpc10*/;
                  if ((13'sd1562/*1562:xpc10*/==xpc10))  xpc10 <= 13'sd1563/*1563:xpc10*/;
                  if ((13'sd1563/*1563:xpc10*/==xpc10))  xpc10 <= 13'sd1564/*1564:xpc10*/;
                  if ((13'sd1565/*1565:xpc10*/==xpc10))  xpc10 <= 13'sd865/*865:xpc10*/;
                  if ((13'sd1566/*1566:xpc10*/==xpc10))  xpc10 <= 13'sd1567/*1567:xpc10*/;
                  if ((13'sd1567/*1567:xpc10*/==xpc10))  xpc10 <= 13'sd1568/*1568:xpc10*/;
                  if ((13'sd1569/*1569:xpc10*/==xpc10))  xpc10 <= 13'sd1562/*1562:xpc10*/;
                  if ((13'sd1570/*1570:xpc10*/==xpc10))  xpc10 <= 13'sd1571/*1571:xpc10*/;
                  if ((13'sd1571/*1571:xpc10*/==xpc10))  xpc10 <= 13'sd1572/*1572:xpc10*/;
                  if ((13'sd1574/*1574:xpc10*/==xpc10))  xpc10 <= 13'sd1081/*1081:xpc10*/;
                  if ((13'sd1575/*1575:xpc10*/==xpc10))  xpc10 <= 13'sd1576/*1576:xpc10*/;
                  if ((13'sd1576/*1576:xpc10*/==xpc10))  xpc10 <= 13'sd1577/*1577:xpc10*/;
                  if ((13'sd1586/*1586:xpc10*/==xpc10))  xpc10 <= 13'sd1587/*1587:xpc10*/;
                  if ((13'sd1587/*1587:xpc10*/==xpc10))  xpc10 <= 13'sd1588/*1588:xpc10*/;
                  if ((13'sd1588/*1588:xpc10*/==xpc10))  xpc10 <= 13'sd1589/*1589:xpc10*/;
                  if ((13'sd1589/*1589:xpc10*/==xpc10))  xpc10 <= 13'sd1590/*1590:xpc10*/;
                  if ((13'sd1590/*1590:xpc10*/==xpc10))  xpc10 <= 13'sd1591/*1591:xpc10*/;
                  if ((13'sd1591/*1591:xpc10*/==xpc10))  xpc10 <= 13'sd1592/*1592:xpc10*/;
                  if ((13'sd1593/*1593:xpc10*/==xpc10))  xpc10 <= 13'sd1594/*1594:xpc10*/;
                  if ((13'sd1594/*1594:xpc10*/==xpc10))  xpc10 <= 13'sd1595/*1595:xpc10*/;
                  if ((13'sd1595/*1595:xpc10*/==xpc10))  xpc10 <= 13'sd1596/*1596:xpc10*/;
                  if ((13'sd1597/*1597:xpc10*/==xpc10))  xpc10 <= 13'sd1598/*1598:xpc10*/;
                  if ((13'sd1598/*1598:xpc10*/==xpc10))  xpc10 <= 13'sd1599/*1599:xpc10*/;
                  if ((13'sd1599/*1599:xpc10*/==xpc10))  xpc10 <= 13'sd1600/*1600:xpc10*/;
                  if ((13'sd1603/*1603:xpc10*/==xpc10))  xpc10 <= 13'sd1604/*1604:xpc10*/;
                  if ((13'sd1604/*1604:xpc10*/==xpc10))  xpc10 <= 13'sd1605/*1605:xpc10*/;
                  if ((13'sd1605/*1605:xpc10*/==xpc10))  xpc10 <= 13'sd1606/*1606:xpc10*/;
                  if ((13'sd1607/*1607:xpc10*/==xpc10))  xpc10 <= 13'sd1608/*1608:xpc10*/;
                  if ((13'sd1608/*1608:xpc10*/==xpc10))  xpc10 <= 13'sd1609/*1609:xpc10*/;
                  if ((13'sd1609/*1609:xpc10*/==xpc10))  xpc10 <= 13'sd1610/*1610:xpc10*/;
                  if ((13'sd1613/*1613:xpc10*/==xpc10))  xpc10 <= 13'sd1614/*1614:xpc10*/;
                  if ((13'sd1614/*1614:xpc10*/==xpc10))  xpc10 <= 13'sd1615/*1615:xpc10*/;
                  if ((13'sd1615/*1615:xpc10*/==xpc10))  xpc10 <= 13'sd1616/*1616:xpc10*/;
                  if ((13'sd1617/*1617:xpc10*/==xpc10))  xpc10 <= 13'sd1618/*1618:xpc10*/;
                  if ((13'sd1618/*1618:xpc10*/==xpc10))  xpc10 <= 13'sd1619/*1619:xpc10*/;
                  if ((13'sd1619/*1619:xpc10*/==xpc10))  xpc10 <= 13'sd1620/*1620:xpc10*/;
                  if ((13'sd1624/*1624:xpc10*/==xpc10))  xpc10 <= 13'sd1625/*1625:xpc10*/;
                  if ((13'sd1625/*1625:xpc10*/==xpc10))  xpc10 <= 13'sd1626/*1626:xpc10*/;
                  if ((13'sd1626/*1626:xpc10*/==xpc10))  xpc10 <= 13'sd1627/*1627:xpc10*/;
                  if ((13'sd1627/*1627:xpc10*/==xpc10))  xpc10 <= 13'sd1628/*1628:xpc10*/;
                  if ((13'sd1628/*1628:xpc10*/==xpc10))  xpc10 <= 13'sd1629/*1629:xpc10*/;
                  if ((13'sd1629/*1629:xpc10*/==xpc10))  xpc10 <= 13'sd1630/*1630:xpc10*/;
                  if ((13'sd1630/*1630:xpc10*/==xpc10))  xpc10 <= 13'sd1631/*1631:xpc10*/;
                  if ((13'sd1632/*1632:xpc10*/==xpc10))  xpc10 <= 13'sd1633/*1633:xpc10*/;
                  if ((13'sd1633/*1633:xpc10*/==xpc10))  xpc10 <= 13'sd1634/*1634:xpc10*/;
                  if ((13'sd1634/*1634:xpc10*/==xpc10))  xpc10 <= 13'sd1635/*1635:xpc10*/;
                  if ((13'sd1636/*1636:xpc10*/==xpc10))  xpc10 <= 13'sd1637/*1637:xpc10*/;
                  if ((13'sd1637/*1637:xpc10*/==xpc10))  xpc10 <= 13'sd1638/*1638:xpc10*/;
                  if ((13'sd1638/*1638:xpc10*/==xpc10))  xpc10 <= 13'sd1639/*1639:xpc10*/;
                  if ((13'sd1640/*1640:xpc10*/==xpc10))  xpc10 <= 13'sd1641/*1641:xpc10*/;
                  if ((13'sd1641/*1641:xpc10*/==xpc10))  xpc10 <= 13'sd1642/*1642:xpc10*/;
                  if ((13'sd1642/*1642:xpc10*/==xpc10))  xpc10 <= 13'sd1643/*1643:xpc10*/;
                  if ((13'sd1644/*1644:xpc10*/==xpc10))  xpc10 <= 13'sd869/*869:xpc10*/;
                  if ((13'sd1645/*1645:xpc10*/==xpc10))  xpc10 <= 13'sd1646/*1646:xpc10*/;
                  if ((13'sd1646/*1646:xpc10*/==xpc10))  xpc10 <= 13'sd1647/*1647:xpc10*/;
                  if ((13'sd1648/*1648:xpc10*/==xpc10))  xpc10 <= 13'sd1649/*1649:xpc10*/;
                  if ((13'sd1649/*1649:xpc10*/==xpc10))  xpc10 <= 13'sd1650/*1650:xpc10*/;
                  if ((13'sd1650/*1650:xpc10*/==xpc10))  xpc10 <= 13'sd1651/*1651:xpc10*/;
                  if ((13'sd1652/*1652:xpc10*/==xpc10))  xpc10 <= 13'sd1637/*1637:xpc10*/;
                  if ((13'sd1653/*1653:xpc10*/==xpc10))  xpc10 <= 13'sd1654/*1654:xpc10*/;
                  if ((13'sd1654/*1654:xpc10*/==xpc10))  xpc10 <= 13'sd1655/*1655:xpc10*/;
                  if ((13'sd1656/*1656:xpc10*/==xpc10))  xpc10 <= 13'sd1657/*1657:xpc10*/;
                  if ((13'sd1657/*1657:xpc10*/==xpc10))  xpc10 <= 13'sd1658/*1658:xpc10*/;
                  if ((13'sd1658/*1658:xpc10*/==xpc10))  xpc10 <= 13'sd1659/*1659:xpc10*/;
                  if ((13'sd1660/*1660:xpc10*/==xpc10))  xpc10 <= 13'sd1637/*1637:xpc10*/;
                  if ((13'sd1661/*1661:xpc10*/==xpc10))  xpc10 <= 13'sd1662/*1662:xpc10*/;
                  if ((13'sd1662/*1662:xpc10*/==xpc10))  xpc10 <= 13'sd1663/*1663:xpc10*/;
                  if ((13'sd1664/*1664:xpc10*/==xpc10))  xpc10 <= 13'sd1637/*1637:xpc10*/;
                  if ((13'sd1665/*1665:xpc10*/==xpc10))  xpc10 <= 13'sd1666/*1666:xpc10*/;
                  if ((13'sd1666/*1666:xpc10*/==xpc10))  xpc10 <= 13'sd1667/*1667:xpc10*/;
                  if ((13'sd1668/*1668:xpc10*/==xpc10))  xpc10 <= 13'sd1618/*1618:xpc10*/;
                  if ((13'sd1669/*1669:xpc10*/==xpc10))  xpc10 <= 13'sd1670/*1670:xpc10*/;
                  if ((13'sd1670/*1670:xpc10*/==xpc10))  xpc10 <= 13'sd1671/*1671:xpc10*/;
                  if ((13'sd1672/*1672:xpc10*/==xpc10))  xpc10 <= 13'sd1608/*1608:xpc10*/;
                  if ((13'sd1673/*1673:xpc10*/==xpc10))  xpc10 <= 13'sd1674/*1674:xpc10*/;
                  if ((13'sd1674/*1674:xpc10*/==xpc10))  xpc10 <= 13'sd1675/*1675:xpc10*/;
                  if ((13'sd1676/*1676:xpc10*/==xpc10))  xpc10 <= 13'sd1641/*1641:xpc10*/;
                  if ((13'sd1677/*1677:xpc10*/==xpc10))  xpc10 <= 13'sd1678/*1678:xpc10*/;
                  if ((13'sd1678/*1678:xpc10*/==xpc10))  xpc10 <= 13'sd1679/*1679:xpc10*/;
                  if ((13'sd1680/*1680:xpc10*/==xpc10))  xpc10 <= 13'sd1681/*1681:xpc10*/;
                  if ((13'sd1681/*1681:xpc10*/==xpc10))  xpc10 <= 13'sd1682/*1682:xpc10*/;
                  if ((13'sd1682/*1682:xpc10*/==xpc10))  xpc10 <= 13'sd1683/*1683:xpc10*/;
                  if ((13'sd1684/*1684:xpc10*/==xpc10))  xpc10 <= 13'sd1685/*1685:xpc10*/;
                  if ((13'sd1685/*1685:xpc10*/==xpc10))  xpc10 <= 13'sd1686/*1686:xpc10*/;
                  if ((13'sd1686/*1686:xpc10*/==xpc10))  xpc10 <= 13'sd1687/*1687:xpc10*/;
                  if ((13'sd1688/*1688:xpc10*/==xpc10))  xpc10 <= 13'sd1689/*1689:xpc10*/;
                  if ((13'sd1689/*1689:xpc10*/==xpc10))  xpc10 <= 13'sd1690/*1690:xpc10*/;
                  if ((13'sd1690/*1690:xpc10*/==xpc10))  xpc10 <= 13'sd1691/*1691:xpc10*/;
                  if ((13'sd1692/*1692:xpc10*/==xpc10))  xpc10 <= 13'sd1693/*1693:xpc10*/;
                  if ((13'sd1693/*1693:xpc10*/==xpc10))  xpc10 <= 13'sd1694/*1694:xpc10*/;
                  if ((13'sd1694/*1694:xpc10*/==xpc10))  xpc10 <= 13'sd1695/*1695:xpc10*/;
                  if ((13'sd1697/*1697:xpc10*/==xpc10))  xpc10 <= 13'sd1698/*1698:xpc10*/;
                  if ((13'sd1698/*1698:xpc10*/==xpc10))  xpc10 <= 13'sd1699/*1699:xpc10*/;
                  if ((13'sd1699/*1699:xpc10*/==xpc10))  xpc10 <= 13'sd1700/*1700:xpc10*/;
                  if ((13'sd1702/*1702:xpc10*/==xpc10))  xpc10 <= 13'sd1703/*1703:xpc10*/;
                  if ((13'sd1703/*1703:xpc10*/==xpc10))  xpc10 <= 13'sd1704/*1704:xpc10*/;
                  if ((13'sd1704/*1704:xpc10*/==xpc10))  xpc10 <= 13'sd1705/*1705:xpc10*/;
                  if ((13'sd1709/*1709:xpc10*/==xpc10))  xpc10 <= 13'sd1710/*1710:xpc10*/;
                  if ((13'sd1710/*1710:xpc10*/==xpc10))  xpc10 <= 13'sd1711/*1711:xpc10*/;
                  if ((13'sd1711/*1711:xpc10*/==xpc10))  xpc10 <= 13'sd1712/*1712:xpc10*/;
                  if ((13'sd1713/*1713:xpc10*/==xpc10))  xpc10 <= 13'sd1714/*1714:xpc10*/;
                  if ((13'sd1714/*1714:xpc10*/==xpc10))  xpc10 <= 13'sd1715/*1715:xpc10*/;
                  if ((13'sd1715/*1715:xpc10*/==xpc10))  xpc10 <= 13'sd1716/*1716:xpc10*/;
                  if ((13'sd1719/*1719:xpc10*/==xpc10))  xpc10 <= 13'sd1720/*1720:xpc10*/;
                  if ((13'sd1720/*1720:xpc10*/==xpc10))  xpc10 <= 13'sd1721/*1721:xpc10*/;
                  if ((13'sd1721/*1721:xpc10*/==xpc10))  xpc10 <= 13'sd1722/*1722:xpc10*/;
                  if ((13'sd1724/*1724:xpc10*/==xpc10))  xpc10 <= 13'sd1725/*1725:xpc10*/;
                  if ((13'sd1725/*1725:xpc10*/==xpc10))  xpc10 <= 13'sd1726/*1726:xpc10*/;
                  if ((13'sd1726/*1726:xpc10*/==xpc10))  xpc10 <= 13'sd1727/*1727:xpc10*/;
                  if ((13'sd1728/*1728:xpc10*/==xpc10))  xpc10 <= 13'sd1729/*1729:xpc10*/;
                  if ((13'sd1729/*1729:xpc10*/==xpc10))  xpc10 <= 13'sd1730/*1730:xpc10*/;
                  if ((13'sd1730/*1730:xpc10*/==xpc10))  xpc10 <= 13'sd1731/*1731:xpc10*/;
                  if ((13'sd1733/*1733:xpc10*/==xpc10))  xpc10 <= 13'sd1734/*1734:xpc10*/;
                  if ((13'sd1734/*1734:xpc10*/==xpc10))  xpc10 <= 13'sd1735/*1735:xpc10*/;
                  if ((13'sd1735/*1735:xpc10*/==xpc10))  xpc10 <= 13'sd1736/*1736:xpc10*/;
                  if ((13'sd1741/*1741:xpc10*/==xpc10))  xpc10 <= 13'sd1742/*1742:xpc10*/;
                  if ((13'sd1742/*1742:xpc10*/==xpc10))  xpc10 <= 13'sd1743/*1743:xpc10*/;
                  if ((13'sd1744/*1744:xpc10*/==xpc10))  xpc10 <= 13'sd1745/*1745:xpc10*/;
                  if ((13'sd1745/*1745:xpc10*/==xpc10))  xpc10 <= 13'sd1746/*1746:xpc10*/;
                  if ((13'sd1746/*1746:xpc10*/==xpc10))  xpc10 <= 13'sd1747/*1747:xpc10*/;
                  if ((13'sd1749/*1749:xpc10*/==xpc10))  xpc10 <= 13'sd1750/*1750:xpc10*/;
                  if ((13'sd1750/*1750:xpc10*/==xpc10))  xpc10 <= 13'sd1751/*1751:xpc10*/;
                  if ((13'sd1751/*1751:xpc10*/==xpc10))  xpc10 <= 13'sd1752/*1752:xpc10*/;
                  if ((13'sd1753/*1753:xpc10*/==xpc10))  xpc10 <= 13'sd1754/*1754:xpc10*/;
                  if ((13'sd1754/*1754:xpc10*/==xpc10))  xpc10 <= 13'sd1755/*1755:xpc10*/;
                  if ((13'sd1755/*1755:xpc10*/==xpc10))  xpc10 <= 13'sd1756/*1756:xpc10*/;
                  if ((13'sd1757/*1757:xpc10*/==xpc10))  xpc10 <= 13'sd1758/*1758:xpc10*/;
                  if ((13'sd1758/*1758:xpc10*/==xpc10))  xpc10 <= 13'sd1759/*1759:xpc10*/;
                  if ((13'sd1759/*1759:xpc10*/==xpc10))  xpc10 <= 13'sd1760/*1760:xpc10*/;
                  if ((13'sd1761/*1761:xpc10*/==xpc10))  xpc10 <= 13'sd1762/*1762:xpc10*/;
                  if ((13'sd1762/*1762:xpc10*/==xpc10))  xpc10 <= 13'sd1763/*1763:xpc10*/;
                  if ((13'sd1763/*1763:xpc10*/==xpc10))  xpc10 <= 13'sd1764/*1764:xpc10*/;
                  if ((13'sd1764/*1764:xpc10*/==xpc10))  xpc10 <= 13'sd1765/*1765:xpc10*/;
                  if ((13'sd1766/*1766:xpc10*/==xpc10))  xpc10 <= 13'sd1767/*1767:xpc10*/;
                  if ((13'sd1767/*1767:xpc10*/==xpc10))  xpc10 <= 13'sd1768/*1768:xpc10*/;
                  if ((13'sd1768/*1768:xpc10*/==xpc10))  xpc10 <= 13'sd1769/*1769:xpc10*/;
                  if ((13'sd1770/*1770:xpc10*/==xpc10))  xpc10 <= 13'sd1771/*1771:xpc10*/;
                  if ((13'sd1771/*1771:xpc10*/==xpc10))  xpc10 <= 13'sd1772/*1772:xpc10*/;
                  if ((13'sd1772/*1772:xpc10*/==xpc10))  xpc10 <= 13'sd1773/*1773:xpc10*/;
                  if ((13'sd1777/*1777:xpc10*/==xpc10))  xpc10 <= 13'sd1778/*1778:xpc10*/;
                  if ((13'sd1778/*1778:xpc10*/==xpc10))  xpc10 <= 13'sd1779/*1779:xpc10*/;
                  if ((13'sd1779/*1779:xpc10*/==xpc10))  xpc10 <= 13'sd1780/*1780:xpc10*/;
                  if ((13'sd1782/*1782:xpc10*/==xpc10))  xpc10 <= 13'sd1783/*1783:xpc10*/;
                  if ((13'sd1783/*1783:xpc10*/==xpc10))  xpc10 <= 13'sd1784/*1784:xpc10*/;
                  if ((13'sd1784/*1784:xpc10*/==xpc10))  xpc10 <= 13'sd1785/*1785:xpc10*/;
                  if ((13'sd1786/*1786:xpc10*/==xpc10))  xpc10 <= 13'sd1787/*1787:xpc10*/;
                  if ((13'sd1787/*1787:xpc10*/==xpc10))  xpc10 <= 13'sd1788/*1788:xpc10*/;
                  if ((13'sd1788/*1788:xpc10*/==xpc10))  xpc10 <= 13'sd1789/*1789:xpc10*/;
                  if ((13'sd1790/*1790:xpc10*/==xpc10))  xpc10 <= 13'sd1641/*1641:xpc10*/;
                  if ((13'sd1791/*1791:xpc10*/==xpc10))  xpc10 <= 13'sd1792/*1792:xpc10*/;
                  if ((13'sd1792/*1792:xpc10*/==xpc10))  xpc10 <= 13'sd1793/*1793:xpc10*/;
                  if ((13'sd1795/*1795:xpc10*/==xpc10))  xpc10 <= 13'sd1783/*1783:xpc10*/;
                  if ((13'sd1796/*1796:xpc10*/==xpc10))  xpc10 <= 13'sd1797/*1797:xpc10*/;
                  if ((13'sd1797/*1797:xpc10*/==xpc10))  xpc10 <= 13'sd1798/*1798:xpc10*/;
                  if ((13'sd1799/*1799:xpc10*/==xpc10))  xpc10 <= 13'sd1771/*1771:xpc10*/;
                  if ((13'sd1800/*1800:xpc10*/==xpc10))  xpc10 <= 13'sd1801/*1801:xpc10*/;
                  if ((13'sd1801/*1801:xpc10*/==xpc10))  xpc10 <= 13'sd1802/*1802:xpc10*/;
                  if ((13'sd1803/*1803:xpc10*/==xpc10))  xpc10 <= 13'sd1804/*1804:xpc10*/;
                  if ((13'sd1804/*1804:xpc10*/==xpc10))  xpc10 <= 13'sd1805/*1805:xpc10*/;
                  if ((13'sd1805/*1805:xpc10*/==xpc10))  xpc10 <= 13'sd1806/*1806:xpc10*/;
                  if ((13'sd1806/*1806:xpc10*/==xpc10))  xpc10 <= 13'sd1807/*1807:xpc10*/;
                  if ((13'sd1808/*1808:xpc10*/==xpc10))  xpc10 <= 13'sd1809/*1809:xpc10*/;
                  if ((13'sd1809/*1809:xpc10*/==xpc10))  xpc10 <= 13'sd1810/*1810:xpc10*/;
                  if ((13'sd1810/*1810:xpc10*/==xpc10))  xpc10 <= 13'sd1811/*1811:xpc10*/;
                  if ((13'sd1812/*1812:xpc10*/==xpc10))  xpc10 <= 13'sd1813/*1813:xpc10*/;
                  if ((13'sd1813/*1813:xpc10*/==xpc10))  xpc10 <= 13'sd1814/*1814:xpc10*/;
                  if ((13'sd1814/*1814:xpc10*/==xpc10))  xpc10 <= 13'sd1815/*1815:xpc10*/;
                  if ((13'sd1818/*1818:xpc10*/==xpc10))  xpc10 <= 13'sd1819/*1819:xpc10*/;
                  if ((13'sd1819/*1819:xpc10*/==xpc10))  xpc10 <= 13'sd1820/*1820:xpc10*/;
                  if ((13'sd1820/*1820:xpc10*/==xpc10))  xpc10 <= 13'sd1821/*1821:xpc10*/;
                  if ((13'sd1822/*1822:xpc10*/==xpc10))  xpc10 <= 13'sd1823/*1823:xpc10*/;
                  if ((13'sd1823/*1823:xpc10*/==xpc10))  xpc10 <= 13'sd1824/*1824:xpc10*/;
                  if ((13'sd1824/*1824:xpc10*/==xpc10))  xpc10 <= 13'sd1825/*1825:xpc10*/;
                  if ((13'sd1825/*1825:xpc10*/==xpc10))  xpc10 <= 13'sd1826/*1826:xpc10*/;
                  if ((13'sd1826/*1826:xpc10*/==xpc10))  xpc10 <= 13'sd1827/*1827:xpc10*/;
                  if ((13'sd1827/*1827:xpc10*/==xpc10))  xpc10 <= 13'sd1828/*1828:xpc10*/;
                  if ((13'sd1828/*1828:xpc10*/==xpc10))  xpc10 <= 13'sd1829/*1829:xpc10*/;
                  if ((13'sd1830/*1830:xpc10*/==xpc10))  xpc10 <= 13'sd1831/*1831:xpc10*/;
                  if ((13'sd1831/*1831:xpc10*/==xpc10))  xpc10 <= 13'sd1832/*1832:xpc10*/;
                  if ((13'sd1832/*1832:xpc10*/==xpc10))  xpc10 <= 13'sd1833/*1833:xpc10*/;
                  if ((13'sd1833/*1833:xpc10*/==xpc10))  xpc10 <= 13'sd1834/*1834:xpc10*/;
                  if ((13'sd1834/*1834:xpc10*/==xpc10))  xpc10 <= 13'sd1835/*1835:xpc10*/;
                  if ((13'sd1835/*1835:xpc10*/==xpc10))  xpc10 <= 13'sd1836/*1836:xpc10*/;
                  if ((13'sd1836/*1836:xpc10*/==xpc10))  xpc10 <= 13'sd1837/*1837:xpc10*/;
                  if ((13'sd1839/*1839:xpc10*/==xpc10))  xpc10 <= 13'sd1840/*1840:xpc10*/;
                  if ((13'sd1840/*1840:xpc10*/==xpc10))  xpc10 <= 13'sd1841/*1841:xpc10*/;
                  if ((13'sd1841/*1841:xpc10*/==xpc10))  xpc10 <= 13'sd1842/*1842:xpc10*/;
                  if ((13'sd1843/*1843:xpc10*/==xpc10))  xpc10 <= 13'sd1844/*1844:xpc10*/;
                  if ((13'sd1844/*1844:xpc10*/==xpc10))  xpc10 <= 13'sd1845/*1845:xpc10*/;
                  if ((13'sd1845/*1845:xpc10*/==xpc10))  xpc10 <= 13'sd1846/*1846:xpc10*/;
                  if ((13'sd1847/*1847:xpc10*/==xpc10))  xpc10 <= 13'sd1848/*1848:xpc10*/;
                  if ((13'sd1848/*1848:xpc10*/==xpc10))  xpc10 <= 13'sd1849/*1849:xpc10*/;
                  if ((13'sd1849/*1849:xpc10*/==xpc10))  xpc10 <= 13'sd1850/*1850:xpc10*/;
                  if ((13'sd1851/*1851:xpc10*/==xpc10))  xpc10 <= 13'sd1852/*1852:xpc10*/;
                  if ((13'sd1852/*1852:xpc10*/==xpc10))  xpc10 <= 13'sd1853/*1853:xpc10*/;
                  if ((13'sd1853/*1853:xpc10*/==xpc10))  xpc10 <= 13'sd1854/*1854:xpc10*/;
                  if ((13'sd1855/*1855:xpc10*/==xpc10))  xpc10 <= 13'sd1856/*1856:xpc10*/;
                  if ((13'sd1856/*1856:xpc10*/==xpc10))  xpc10 <= 13'sd1857/*1857:xpc10*/;
                  if ((13'sd1857/*1857:xpc10*/==xpc10))  xpc10 <= 13'sd1858/*1858:xpc10*/;
                  if ((13'sd1859/*1859:xpc10*/==xpc10))  xpc10 <= 13'sd1860/*1860:xpc10*/;
                  if ((13'sd1860/*1860:xpc10*/==xpc10))  xpc10 <= 13'sd1861/*1861:xpc10*/;
                  if ((13'sd1861/*1861:xpc10*/==xpc10))  xpc10 <= 13'sd1862/*1862:xpc10*/;
                  if ((13'sd1863/*1863:xpc10*/==xpc10))  xpc10 <= 13'sd1787/*1787:xpc10*/;
                  if ((13'sd1864/*1864:xpc10*/==xpc10))  xpc10 <= 13'sd1865/*1865:xpc10*/;
                  if ((13'sd1865/*1865:xpc10*/==xpc10))  xpc10 <= 13'sd1866/*1866:xpc10*/;
                  if ((13'sd1867/*1867:xpc10*/==xpc10))  xpc10 <= 13'sd1860/*1860:xpc10*/;
                  if ((13'sd1868/*1868:xpc10*/==xpc10))  xpc10 <= 13'sd1869/*1869:xpc10*/;
                  if ((13'sd1869/*1869:xpc10*/==xpc10))  xpc10 <= 13'sd1870/*1870:xpc10*/;
                  if ((13'sd1871/*1871:xpc10*/==xpc10))  xpc10 <= 13'sd1872/*1872:xpc10*/;
                  if ((13'sd1872/*1872:xpc10*/==xpc10))  xpc10 <= 13'sd1873/*1873:xpc10*/;
                  if ((13'sd1873/*1873:xpc10*/==xpc10))  xpc10 <= 13'sd1874/*1874:xpc10*/;
                  if ((13'sd1878/*1878:xpc10*/==xpc10))  xpc10 <= 13'sd1879/*1879:xpc10*/;
                  if ((13'sd1879/*1879:xpc10*/==xpc10))  xpc10 <= 13'sd1880/*1880:xpc10*/;
                  if ((13'sd1880/*1880:xpc10*/==xpc10))  xpc10 <= 13'sd1881/*1881:xpc10*/;
                  if ((13'sd1883/*1883:xpc10*/==xpc10))  xpc10 <= 13'sd1884/*1884:xpc10*/;
                  if ((13'sd1884/*1884:xpc10*/==xpc10))  xpc10 <= 13'sd1885/*1885:xpc10*/;
                  if ((13'sd1885/*1885:xpc10*/==xpc10))  xpc10 <= 13'sd1886/*1886:xpc10*/;
                  if ((13'sd1887/*1887:xpc10*/==xpc10))  xpc10 <= 13'sd1813/*1813:xpc10*/;
                  if ((13'sd1888/*1888:xpc10*/==xpc10))  xpc10 <= 13'sd1889/*1889:xpc10*/;
                  if ((13'sd1889/*1889:xpc10*/==xpc10))  xpc10 <= 13'sd1890/*1890:xpc10*/;
                  if ((13'sd1892/*1892:xpc10*/==xpc10))  xpc10 <= 13'sd1884/*1884:xpc10*/;
                  if ((13'sd1893/*1893:xpc10*/==xpc10))  xpc10 <= 13'sd1894/*1894:xpc10*/;
                  if ((13'sd1894/*1894:xpc10*/==xpc10))  xpc10 <= 13'sd1895/*1895:xpc10*/;
                  if ((13'sd1896/*1896:xpc10*/==xpc10))  xpc10 <= 13'sd1897/*1897:xpc10*/;
                  if ((13'sd1897/*1897:xpc10*/==xpc10))  xpc10 <= 13'sd1898/*1898:xpc10*/;
                  if ((13'sd1898/*1898:xpc10*/==xpc10))  xpc10 <= 13'sd1899/*1899:xpc10*/;
                  if ((13'sd1900/*1900:xpc10*/==xpc10))  xpc10 <= 13'sd1901/*1901:xpc10*/;
                  if ((13'sd1901/*1901:xpc10*/==xpc10))  xpc10 <= 13'sd1902/*1902:xpc10*/;
                  if ((13'sd1902/*1902:xpc10*/==xpc10))  xpc10 <= 13'sd1903/*1903:xpc10*/;
                  if ((13'sd1904/*1904:xpc10*/==xpc10))  xpc10 <= 13'sd1813/*1813:xpc10*/;
                  if ((13'sd1905/*1905:xpc10*/==xpc10))  xpc10 <= 13'sd1906/*1906:xpc10*/;
                  if ((13'sd1906/*1906:xpc10*/==xpc10))  xpc10 <= 13'sd1907/*1907:xpc10*/;
                  if ((13'sd1908/*1908:xpc10*/==xpc10))  xpc10 <= 13'sd1901/*1901:xpc10*/;
                  if ((13'sd1909/*1909:xpc10*/==xpc10))  xpc10 <= 13'sd1910/*1910:xpc10*/;
                  if ((13'sd1910/*1910:xpc10*/==xpc10))  xpc10 <= 13'sd1911/*1911:xpc10*/;
                  if ((13'sd1912/*1912:xpc10*/==xpc10))  xpc10 <= 13'sd1714/*1714:xpc10*/;
                  if ((13'sd1913/*1913:xpc10*/==xpc10))  xpc10 <= 13'sd1914/*1914:xpc10*/;
                  if ((13'sd1914/*1914:xpc10*/==xpc10))  xpc10 <= 13'sd1915/*1915:xpc10*/;
                  if ((13'sd1916/*1916:xpc10*/==xpc10))  xpc10 <= 13'sd1917/*1917:xpc10*/;
                  if ((13'sd1917/*1917:xpc10*/==xpc10))  xpc10 <= 13'sd1918/*1918:xpc10*/;
                  if ((13'sd1918/*1918:xpc10*/==xpc10))  xpc10 <= 13'sd1919/*1919:xpc10*/;
                  if ((13'sd1923/*1923:xpc10*/==xpc10))  xpc10 <= 13'sd1924/*1924:xpc10*/;
                  if ((13'sd1924/*1924:xpc10*/==xpc10))  xpc10 <= 13'sd1925/*1925:xpc10*/;
                  if ((13'sd1925/*1925:xpc10*/==xpc10))  xpc10 <= 13'sd1926/*1926:xpc10*/;
                  if ((13'sd1928/*1928:xpc10*/==xpc10))  xpc10 <= 13'sd1929/*1929:xpc10*/;
                  if ((13'sd1929/*1929:xpc10*/==xpc10))  xpc10 <= 13'sd1930/*1930:xpc10*/;
                  if ((13'sd1930/*1930:xpc10*/==xpc10))  xpc10 <= 13'sd1931/*1931:xpc10*/;
                  if ((13'sd1932/*1932:xpc10*/==xpc10))  xpc10 <= 13'sd1693/*1693:xpc10*/;
                  if ((13'sd1933/*1933:xpc10*/==xpc10))  xpc10 <= 13'sd1934/*1934:xpc10*/;
                  if ((13'sd1934/*1934:xpc10*/==xpc10))  xpc10 <= 13'sd1935/*1935:xpc10*/;
                  if ((13'sd1937/*1937:xpc10*/==xpc10))  xpc10 <= 13'sd1929/*1929:xpc10*/;
                  if ((13'sd1938/*1938:xpc10*/==xpc10))  xpc10 <= 13'sd1939/*1939:xpc10*/;
                  if ((13'sd1939/*1939:xpc10*/==xpc10))  xpc10 <= 13'sd1940/*1940:xpc10*/;
                  if ((13'sd1941/*1941:xpc10*/==xpc10))  xpc10 <= 13'sd1942/*1942:xpc10*/;
                  if ((13'sd1942/*1942:xpc10*/==xpc10))  xpc10 <= 13'sd1943/*1943:xpc10*/;
                  if ((13'sd1943/*1943:xpc10*/==xpc10))  xpc10 <= 13'sd1944/*1944:xpc10*/;
                  if ((13'sd1945/*1945:xpc10*/==xpc10))  xpc10 <= 13'sd1946/*1946:xpc10*/;
                  if ((13'sd1946/*1946:xpc10*/==xpc10))  xpc10 <= 13'sd1947/*1947:xpc10*/;
                  if ((13'sd1947/*1947:xpc10*/==xpc10))  xpc10 <= 13'sd1948/*1948:xpc10*/;
                  if ((13'sd1949/*1949:xpc10*/==xpc10))  xpc10 <= 13'sd1693/*1693:xpc10*/;
                  if ((13'sd1950/*1950:xpc10*/==xpc10))  xpc10 <= 13'sd1951/*1951:xpc10*/;
                  if ((13'sd1951/*1951:xpc10*/==xpc10))  xpc10 <= 13'sd1952/*1952:xpc10*/;
                  if ((13'sd1953/*1953:xpc10*/==xpc10))  xpc10 <= 13'sd1946/*1946:xpc10*/;
                  if ((13'sd1954/*1954:xpc10*/==xpc10))  xpc10 <= 13'sd1955/*1955:xpc10*/;
                  if ((13'sd1955/*1955:xpc10*/==xpc10))  xpc10 <= 13'sd1956/*1956:xpc10*/;
                  if ((13'sd1957/*1957:xpc10*/==xpc10))  xpc10 <= 13'sd1685/*1685:xpc10*/;
                  if ((13'sd1958/*1958:xpc10*/==xpc10))  xpc10 <= 13'sd1959/*1959:xpc10*/;
                  if ((13'sd1959/*1959:xpc10*/==xpc10))  xpc10 <= 13'sd1960/*1960:xpc10*/;
                  if ((13'sd1961/*1961:xpc10*/==xpc10))  xpc10 <= 13'sd1962/*1962:xpc10*/;
                  if ((13'sd1962/*1962:xpc10*/==xpc10))  xpc10 <= 13'sd1963/*1963:xpc10*/;
                  if ((13'sd1963/*1963:xpc10*/==xpc10))  xpc10 <= 13'sd1964/*1964:xpc10*/;
                  if ((13'sd1964/*1964:xpc10*/==xpc10))  xpc10 <= 13'sd1965/*1965:xpc10*/;
                  if ((13'sd1965/*1965:xpc10*/==xpc10))  xpc10 <= 13'sd1966/*1966:xpc10*/;
                  if ((13'sd1966/*1966:xpc10*/==xpc10))  xpc10 <= 13'sd1967/*1967:xpc10*/;
                  if ((13'sd1968/*1968:xpc10*/==xpc10))  xpc10 <= 13'sd1969/*1969:xpc10*/;
                  if ((13'sd1969/*1969:xpc10*/==xpc10))  xpc10 <= 13'sd1970/*1970:xpc10*/;
                  if ((13'sd1970/*1970:xpc10*/==xpc10))  xpc10 <= 13'sd1971/*1971:xpc10*/;
                  if ((13'sd1972/*1972:xpc10*/==xpc10))  xpc10 <= 13'sd1973/*1973:xpc10*/;
                  if ((13'sd1973/*1973:xpc10*/==xpc10))  xpc10 <= 13'sd1974/*1974:xpc10*/;
                  if ((13'sd1974/*1974:xpc10*/==xpc10))  xpc10 <= 13'sd1975/*1975:xpc10*/;
                  if ((13'sd1978/*1978:xpc10*/==xpc10))  xpc10 <= 13'sd1979/*1979:xpc10*/;
                  if ((13'sd1979/*1979:xpc10*/==xpc10))  xpc10 <= 13'sd1980/*1980:xpc10*/;
                  if ((13'sd1980/*1980:xpc10*/==xpc10))  xpc10 <= 13'sd1981/*1981:xpc10*/;
                  if ((13'sd1982/*1982:xpc10*/==xpc10))  xpc10 <= 13'sd1983/*1983:xpc10*/;
                  if ((13'sd1983/*1983:xpc10*/==xpc10))  xpc10 <= 13'sd1984/*1984:xpc10*/;
                  if ((13'sd1984/*1984:xpc10*/==xpc10))  xpc10 <= 13'sd1985/*1985:xpc10*/;
                  if ((13'sd1988/*1988:xpc10*/==xpc10))  xpc10 <= 13'sd1989/*1989:xpc10*/;
                  if ((13'sd1989/*1989:xpc10*/==xpc10))  xpc10 <= 13'sd1990/*1990:xpc10*/;
                  if ((13'sd1990/*1990:xpc10*/==xpc10))  xpc10 <= 13'sd1991/*1991:xpc10*/;
                  if ((13'sd1992/*1992:xpc10*/==xpc10))  xpc10 <= 13'sd1993/*1993:xpc10*/;
                  if ((13'sd1993/*1993:xpc10*/==xpc10))  xpc10 <= 13'sd1994/*1994:xpc10*/;
                  if ((13'sd1994/*1994:xpc10*/==xpc10))  xpc10 <= 13'sd1995/*1995:xpc10*/;
                  if ((13'sd1999/*1999:xpc10*/==xpc10))  xpc10 <= 13'sd2000/*2000:xpc10*/;
                  if ((13'sd2000/*2000:xpc10*/==xpc10))  xpc10 <= 13'sd2001/*2001:xpc10*/;
                  if ((13'sd2001/*2001:xpc10*/==xpc10))  xpc10 <= 13'sd2002/*2002:xpc10*/;
                  if ((13'sd2002/*2002:xpc10*/==xpc10))  xpc10 <= 13'sd2003/*2003:xpc10*/;
                  if ((13'sd2003/*2003:xpc10*/==xpc10))  xpc10 <= 13'sd2004/*2004:xpc10*/;
                  if ((13'sd2004/*2004:xpc10*/==xpc10))  xpc10 <= 13'sd2005/*2005:xpc10*/;
                  if ((13'sd2005/*2005:xpc10*/==xpc10))  xpc10 <= 13'sd2006/*2006:xpc10*/;
                  if ((13'sd2007/*2007:xpc10*/==xpc10))  xpc10 <= 13'sd2008/*2008:xpc10*/;
                  if ((13'sd2008/*2008:xpc10*/==xpc10))  xpc10 <= 13'sd2009/*2009:xpc10*/;
                  if ((13'sd2009/*2009:xpc10*/==xpc10))  xpc10 <= 13'sd2010/*2010:xpc10*/;
                  if ((13'sd2011/*2011:xpc10*/==xpc10))  xpc10 <= 13'sd2012/*2012:xpc10*/;
                  if ((13'sd2012/*2012:xpc10*/==xpc10))  xpc10 <= 13'sd2013/*2013:xpc10*/;
                  if ((13'sd2013/*2013:xpc10*/==xpc10))  xpc10 <= 13'sd2014/*2014:xpc10*/;
                  if ((13'sd2015/*2015:xpc10*/==xpc10))  xpc10 <= 13'sd1641/*1641:xpc10*/;
                  if ((13'sd2016/*2016:xpc10*/==xpc10))  xpc10 <= 13'sd2017/*2017:xpc10*/;
                  if ((13'sd2017/*2017:xpc10*/==xpc10))  xpc10 <= 13'sd2018/*2018:xpc10*/;
                  if ((13'sd2019/*2019:xpc10*/==xpc10))  xpc10 <= 13'sd2020/*2020:xpc10*/;
                  if ((13'sd2020/*2020:xpc10*/==xpc10))  xpc10 <= 13'sd2021/*2021:xpc10*/;
                  if ((13'sd2021/*2021:xpc10*/==xpc10))  xpc10 <= 13'sd2022/*2022:xpc10*/;
                  if ((13'sd2023/*2023:xpc10*/==xpc10))  xpc10 <= 13'sd2012/*2012:xpc10*/;
                  if ((13'sd2024/*2024:xpc10*/==xpc10))  xpc10 <= 13'sd2025/*2025:xpc10*/;
                  if ((13'sd2025/*2025:xpc10*/==xpc10))  xpc10 <= 13'sd2026/*2026:xpc10*/;
                  if ((13'sd2027/*2027:xpc10*/==xpc10))  xpc10 <= 13'sd2028/*2028:xpc10*/;
                  if ((13'sd2028/*2028:xpc10*/==xpc10))  xpc10 <= 13'sd2029/*2029:xpc10*/;
                  if ((13'sd2029/*2029:xpc10*/==xpc10))  xpc10 <= 13'sd2030/*2030:xpc10*/;
                  if ((13'sd2031/*2031:xpc10*/==xpc10))  xpc10 <= 13'sd2012/*2012:xpc10*/;
                  if ((13'sd2032/*2032:xpc10*/==xpc10))  xpc10 <= 13'sd2033/*2033:xpc10*/;
                  if ((13'sd2033/*2033:xpc10*/==xpc10))  xpc10 <= 13'sd2034/*2034:xpc10*/;
                  if ((13'sd2035/*2035:xpc10*/==xpc10))  xpc10 <= 13'sd2012/*2012:xpc10*/;
                  if ((13'sd2036/*2036:xpc10*/==xpc10))  xpc10 <= 13'sd2037/*2037:xpc10*/;
                  if ((13'sd2037/*2037:xpc10*/==xpc10))  xpc10 <= 13'sd2038/*2038:xpc10*/;
                  if ((13'sd2039/*2039:xpc10*/==xpc10))  xpc10 <= 13'sd1993/*1993:xpc10*/;
                  if ((13'sd2040/*2040:xpc10*/==xpc10))  xpc10 <= 13'sd2041/*2041:xpc10*/;
                  if ((13'sd2041/*2041:xpc10*/==xpc10))  xpc10 <= 13'sd2042/*2042:xpc10*/;
                  if ((13'sd2043/*2043:xpc10*/==xpc10))  xpc10 <= 13'sd1983/*1983:xpc10*/;
                  if ((13'sd2044/*2044:xpc10*/==xpc10))  xpc10 <= 13'sd2045/*2045:xpc10*/;
                  if ((13'sd2045/*2045:xpc10*/==xpc10))  xpc10 <= 13'sd2046/*2046:xpc10*/;
                  if ((13'sd2047/*2047:xpc10*/==xpc10))  xpc10 <= 13'sd2048/*2048:xpc10*/;
                  if ((13'sd2048/*2048:xpc10*/==xpc10))  xpc10 <= 13'sd2049/*2049:xpc10*/;
                  if ((13'sd2049/*2049:xpc10*/==xpc10))  xpc10 <= 13'sd2050/*2050:xpc10*/;
                  if ((13'sd2051/*2051:xpc10*/==xpc10))  xpc10 <= 13'sd2052/*2052:xpc10*/;
                  if ((13'sd2052/*2052:xpc10*/==xpc10))  xpc10 <= 13'sd2053/*2053:xpc10*/;
                  if ((13'sd2053/*2053:xpc10*/==xpc10))  xpc10 <= 13'sd2054/*2054:xpc10*/;
                  if ((13'sd2055/*2055:xpc10*/==xpc10))  xpc10 <= 13'sd1641/*1641:xpc10*/;
                  if ((13'sd2056/*2056:xpc10*/==xpc10))  xpc10 <= 13'sd2057/*2057:xpc10*/;
                  if ((13'sd2057/*2057:xpc10*/==xpc10))  xpc10 <= 13'sd2058/*2058:xpc10*/;
                  if ((13'sd2059/*2059:xpc10*/==xpc10))  xpc10 <= 13'sd2052/*2052:xpc10*/;
                  if ((13'sd2060/*2060:xpc10*/==xpc10))  xpc10 <= 13'sd2061/*2061:xpc10*/;
                  if ((13'sd2061/*2061:xpc10*/==xpc10))  xpc10 <= 13'sd2062/*2062:xpc10*/;
                  if ((13'sd2063/*2063:xpc10*/==xpc10))  xpc10 <= 13'sd2064/*2064:xpc10*/;
                  if ((13'sd2064/*2064:xpc10*/==xpc10))  xpc10 <= 13'sd2065/*2065:xpc10*/;
                  if ((13'sd2065/*2065:xpc10*/==xpc10))  xpc10 <= 13'sd2066/*2066:xpc10*/;
                  if ((13'sd2067/*2067:xpc10*/==xpc10))  xpc10 <= 13'sd2068/*2068:xpc10*/;
                  if ((13'sd2068/*2068:xpc10*/==xpc10))  xpc10 <= 13'sd2069/*2069:xpc10*/;
                  if ((13'sd2069/*2069:xpc10*/==xpc10))  xpc10 <= 13'sd2070/*2070:xpc10*/;
                  if ((13'sd2071/*2071:xpc10*/==xpc10))  xpc10 <= 13'sd2072/*2072:xpc10*/;
                  if ((13'sd2072/*2072:xpc10*/==xpc10))  xpc10 <= 13'sd2073/*2073:xpc10*/;
                  if ((13'sd2073/*2073:xpc10*/==xpc10))  xpc10 <= 13'sd2074/*2074:xpc10*/;
                  if ((13'sd2075/*2075:xpc10*/==xpc10))  xpc10 <= 13'sd2076/*2076:xpc10*/;
                  if ((13'sd2076/*2076:xpc10*/==xpc10))  xpc10 <= 13'sd2077/*2077:xpc10*/;
                  if ((13'sd2077/*2077:xpc10*/==xpc10))  xpc10 <= 13'sd2078/*2078:xpc10*/;
                  if ((13'sd2080/*2080:xpc10*/==xpc10))  xpc10 <= 13'sd2081/*2081:xpc10*/;
                  if ((13'sd2081/*2081:xpc10*/==xpc10))  xpc10 <= 13'sd2082/*2082:xpc10*/;
                  if ((13'sd2082/*2082:xpc10*/==xpc10))  xpc10 <= 13'sd2083/*2083:xpc10*/;
                  if ((13'sd2086/*2086:xpc10*/==xpc10))  xpc10 <= 13'sd1703/*1703:xpc10*/;
                  if ((13'sd2087/*2087:xpc10*/==xpc10))  xpc10 <= 13'sd2088/*2088:xpc10*/;
                  if ((13'sd2088/*2088:xpc10*/==xpc10))  xpc10 <= 13'sd2089/*2089:xpc10*/;
                  if ((13'sd2090/*2090:xpc10*/==xpc10))  xpc10 <= 13'sd2091/*2091:xpc10*/;
                  if ((13'sd2091/*2091:xpc10*/==xpc10))  xpc10 <= 13'sd2092/*2092:xpc10*/;
                  if ((13'sd2092/*2092:xpc10*/==xpc10))  xpc10 <= 13'sd2093/*2093:xpc10*/;
                  if ((13'sd2097/*2097:xpc10*/==xpc10))  xpc10 <= 13'sd2098/*2098:xpc10*/;
                  if ((13'sd2098/*2098:xpc10*/==xpc10))  xpc10 <= 13'sd2099/*2099:xpc10*/;
                  if ((13'sd2099/*2099:xpc10*/==xpc10))  xpc10 <= 13'sd2100/*2100:xpc10*/;
                  if ((13'sd2102/*2102:xpc10*/==xpc10))  xpc10 <= 13'sd2103/*2103:xpc10*/;
                  if ((13'sd2103/*2103:xpc10*/==xpc10))  xpc10 <= 13'sd2104/*2104:xpc10*/;
                  if ((13'sd2104/*2104:xpc10*/==xpc10))  xpc10 <= 13'sd2105/*2105:xpc10*/;
                  if ((13'sd2106/*2106:xpc10*/==xpc10))  xpc10 <= 13'sd2076/*2076:xpc10*/;
                  if ((13'sd2107/*2107:xpc10*/==xpc10))  xpc10 <= 13'sd2108/*2108:xpc10*/;
                  if ((13'sd2108/*2108:xpc10*/==xpc10))  xpc10 <= 13'sd2109/*2109:xpc10*/;
                  if ((13'sd2111/*2111:xpc10*/==xpc10))  xpc10 <= 13'sd2103/*2103:xpc10*/;
                  if ((13'sd2112/*2112:xpc10*/==xpc10))  xpc10 <= 13'sd2113/*2113:xpc10*/;
                  if ((13'sd2113/*2113:xpc10*/==xpc10))  xpc10 <= 13'sd2114/*2114:xpc10*/;
                  if ((13'sd2115/*2115:xpc10*/==xpc10))  xpc10 <= 13'sd2116/*2116:xpc10*/;
                  if ((13'sd2116/*2116:xpc10*/==xpc10))  xpc10 <= 13'sd2117/*2117:xpc10*/;
                  if ((13'sd2117/*2117:xpc10*/==xpc10))  xpc10 <= 13'sd2118/*2118:xpc10*/;
                  if ((13'sd2119/*2119:xpc10*/==xpc10))  xpc10 <= 13'sd2120/*2120:xpc10*/;
                  if ((13'sd2120/*2120:xpc10*/==xpc10))  xpc10 <= 13'sd2121/*2121:xpc10*/;
                  if ((13'sd2121/*2121:xpc10*/==xpc10))  xpc10 <= 13'sd2122/*2122:xpc10*/;
                  if ((13'sd2123/*2123:xpc10*/==xpc10))  xpc10 <= 13'sd2076/*2076:xpc10*/;
                  if ((13'sd2124/*2124:xpc10*/==xpc10))  xpc10 <= 13'sd2125/*2125:xpc10*/;
                  if ((13'sd2125/*2125:xpc10*/==xpc10))  xpc10 <= 13'sd2126/*2126:xpc10*/;
                  if ((13'sd2127/*2127:xpc10*/==xpc10))  xpc10 <= 13'sd2120/*2120:xpc10*/;
                  if ((13'sd2128/*2128:xpc10*/==xpc10))  xpc10 <= 13'sd2129/*2129:xpc10*/;
                  if ((13'sd2129/*2129:xpc10*/==xpc10))  xpc10 <= 13'sd2130/*2130:xpc10*/;
                  if ((13'sd2131/*2131:xpc10*/==xpc10))  xpc10 <= 13'sd2068/*2068:xpc10*/;
                  if ((13'sd2132/*2132:xpc10*/==xpc10))  xpc10 <= 13'sd2133/*2133:xpc10*/;
                  if ((13'sd2133/*2133:xpc10*/==xpc10))  xpc10 <= 13'sd2134/*2134:xpc10*/;
                  if ((13'sd2135/*2135:xpc10*/==xpc10))  xpc10 <= 13'sd2136/*2136:xpc10*/;
                  if ((13'sd2136/*2136:xpc10*/==xpc10))  xpc10 <= 13'sd2137/*2137:xpc10*/;
                  if ((13'sd2137/*2137:xpc10*/==xpc10))  xpc10 <= 13'sd2138/*2138:xpc10*/;
                  if ((13'sd2139/*2139:xpc10*/==xpc10))  xpc10 <= 13'sd2140/*2140:xpc10*/;
                  if ((13'sd2140/*2140:xpc10*/==xpc10))  xpc10 <= 13'sd2141/*2141:xpc10*/;
                  if ((13'sd2141/*2141:xpc10*/==xpc10))  xpc10 <= 13'sd2142/*2142:xpc10*/;
                  if ((13'sd2143/*2143:xpc10*/==xpc10))  xpc10 <= 13'sd2144/*2144:xpc10*/;
                  if ((13'sd2144/*2144:xpc10*/==xpc10))  xpc10 <= 13'sd2145/*2145:xpc10*/;
                  if ((13'sd2145/*2145:xpc10*/==xpc10))  xpc10 <= 13'sd2146/*2146:xpc10*/;
                  if ((13'sd2149/*2149:xpc10*/==xpc10))  xpc10 <= 13'sd2150/*2150:xpc10*/;
                  if ((13'sd2150/*2150:xpc10*/==xpc10))  xpc10 <= 13'sd2151/*2151:xpc10*/;
                  if ((13'sd2151/*2151:xpc10*/==xpc10))  xpc10 <= 13'sd2152/*2152:xpc10*/;
                  if ((13'sd2153/*2153:xpc10*/==xpc10))  xpc10 <= 13'sd2154/*2154:xpc10*/;
                  if ((13'sd2154/*2154:xpc10*/==xpc10))  xpc10 <= 13'sd2155/*2155:xpc10*/;
                  if ((13'sd2155/*2155:xpc10*/==xpc10))  xpc10 <= 13'sd2156/*2156:xpc10*/;
                  if ((13'sd2159/*2159:xpc10*/==xpc10))  xpc10 <= 13'sd2160/*2160:xpc10*/;
                  if ((13'sd2160/*2160:xpc10*/==xpc10))  xpc10 <= 13'sd2161/*2161:xpc10*/;
                  if ((13'sd2161/*2161:xpc10*/==xpc10))  xpc10 <= 13'sd2162/*2162:xpc10*/;
                  if ((13'sd2163/*2163:xpc10*/==xpc10))  xpc10 <= 13'sd2164/*2164:xpc10*/;
                  if ((13'sd2164/*2164:xpc10*/==xpc10))  xpc10 <= 13'sd2165/*2165:xpc10*/;
                  if ((13'sd2165/*2165:xpc10*/==xpc10))  xpc10 <= 13'sd2166/*2166:xpc10*/;
                  if ((13'sd2170/*2170:xpc10*/==xpc10))  xpc10 <= 13'sd2171/*2171:xpc10*/;
                  if ((13'sd2171/*2171:xpc10*/==xpc10))  xpc10 <= 13'sd2172/*2172:xpc10*/;
                  if ((13'sd2172/*2172:xpc10*/==xpc10))  xpc10 <= 13'sd2173/*2173:xpc10*/;
                  if ((13'sd2173/*2173:xpc10*/==xpc10))  xpc10 <= 13'sd2174/*2174:xpc10*/;
                  if ((13'sd2174/*2174:xpc10*/==xpc10))  xpc10 <= 13'sd2175/*2175:xpc10*/;
                  if ((13'sd2175/*2175:xpc10*/==xpc10))  xpc10 <= 13'sd2176/*2176:xpc10*/;
                  if ((13'sd2176/*2176:xpc10*/==xpc10))  xpc10 <= 13'sd2177/*2177:xpc10*/;
                  if ((13'sd2178/*2178:xpc10*/==xpc10))  xpc10 <= 13'sd2179/*2179:xpc10*/;
                  if ((13'sd2179/*2179:xpc10*/==xpc10))  xpc10 <= 13'sd2180/*2180:xpc10*/;
                  if ((13'sd2180/*2180:xpc10*/==xpc10))  xpc10 <= 13'sd2181/*2181:xpc10*/;
                  if ((13'sd2182/*2182:xpc10*/==xpc10))  xpc10 <= 13'sd2183/*2183:xpc10*/;
                  if ((13'sd2183/*2183:xpc10*/==xpc10))  xpc10 <= 13'sd2184/*2184:xpc10*/;
                  if ((13'sd2184/*2184:xpc10*/==xpc10))  xpc10 <= 13'sd2185/*2185:xpc10*/;
                  if ((13'sd2186/*2186:xpc10*/==xpc10))  xpc10 <= 13'sd1641/*1641:xpc10*/;
                  if ((13'sd2187/*2187:xpc10*/==xpc10))  xpc10 <= 13'sd2188/*2188:xpc10*/;
                  if ((13'sd2188/*2188:xpc10*/==xpc10))  xpc10 <= 13'sd2189/*2189:xpc10*/;
                  if ((13'sd2190/*2190:xpc10*/==xpc10))  xpc10 <= 13'sd2191/*2191:xpc10*/;
                  if ((13'sd2191/*2191:xpc10*/==xpc10))  xpc10 <= 13'sd2192/*2192:xpc10*/;
                  if ((13'sd2192/*2192:xpc10*/==xpc10))  xpc10 <= 13'sd2193/*2193:xpc10*/;
                  if ((13'sd2194/*2194:xpc10*/==xpc10))  xpc10 <= 13'sd2183/*2183:xpc10*/;
                  if ((13'sd2195/*2195:xpc10*/==xpc10))  xpc10 <= 13'sd2196/*2196:xpc10*/;
                  if ((13'sd2196/*2196:xpc10*/==xpc10))  xpc10 <= 13'sd2197/*2197:xpc10*/;
                  if ((13'sd2198/*2198:xpc10*/==xpc10))  xpc10 <= 13'sd2199/*2199:xpc10*/;
                  if ((13'sd2199/*2199:xpc10*/==xpc10))  xpc10 <= 13'sd2200/*2200:xpc10*/;
                  if ((13'sd2200/*2200:xpc10*/==xpc10))  xpc10 <= 13'sd2201/*2201:xpc10*/;
                  if ((13'sd2202/*2202:xpc10*/==xpc10))  xpc10 <= 13'sd2183/*2183:xpc10*/;
                  if ((13'sd2203/*2203:xpc10*/==xpc10))  xpc10 <= 13'sd2204/*2204:xpc10*/;
                  if ((13'sd2204/*2204:xpc10*/==xpc10))  xpc10 <= 13'sd2205/*2205:xpc10*/;
                  if ((13'sd2206/*2206:xpc10*/==xpc10))  xpc10 <= 13'sd2183/*2183:xpc10*/;
                  if ((13'sd2207/*2207:xpc10*/==xpc10))  xpc10 <= 13'sd2208/*2208:xpc10*/;
                  if ((13'sd2208/*2208:xpc10*/==xpc10))  xpc10 <= 13'sd2209/*2209:xpc10*/;
                  if ((13'sd2210/*2210:xpc10*/==xpc10))  xpc10 <= 13'sd2164/*2164:xpc10*/;
                  if ((13'sd2211/*2211:xpc10*/==xpc10))  xpc10 <= 13'sd2212/*2212:xpc10*/;
                  if ((13'sd2212/*2212:xpc10*/==xpc10))  xpc10 <= 13'sd2213/*2213:xpc10*/;
                  if ((13'sd2214/*2214:xpc10*/==xpc10))  xpc10 <= 13'sd2154/*2154:xpc10*/;
                  if ((13'sd2215/*2215:xpc10*/==xpc10))  xpc10 <= 13'sd2216/*2216:xpc10*/;
                  if ((13'sd2216/*2216:xpc10*/==xpc10))  xpc10 <= 13'sd2217/*2217:xpc10*/;
                  if ((13'sd2217/*2217:xpc10*/==xpc10))  xpc10 <= 13'sd2218/*2218:xpc10*/;
                  if ((13'sd2219/*2219:xpc10*/==xpc10))  xpc10 <= 13'sd1641/*1641:xpc10*/;
                  if ((13'sd2220/*2220:xpc10*/==xpc10))  xpc10 <= 13'sd2221/*2221:xpc10*/;
                  if ((13'sd2221/*2221:xpc10*/==xpc10))  xpc10 <= 13'sd2222/*2222:xpc10*/;
                  if ((13'sd2223/*2223:xpc10*/==xpc10))  xpc10 <= 13'sd2224/*2224:xpc10*/;
                  if ((13'sd2224/*2224:xpc10*/==xpc10))  xpc10 <= 13'sd2225/*2225:xpc10*/;
                  if ((13'sd2225/*2225:xpc10*/==xpc10))  xpc10 <= 13'sd2226/*2226:xpc10*/;
                  if ((13'sd2228/*2228:xpc10*/==xpc10))  xpc10 <= 13'sd2229/*2229:xpc10*/;
                  if ((13'sd2229/*2229:xpc10*/==xpc10))  xpc10 <= 13'sd2230/*2230:xpc10*/;
                  if ((13'sd2230/*2230:xpc10*/==xpc10))  xpc10 <= 13'sd2231/*2231:xpc10*/;
                  if ((13'sd2232/*2232:xpc10*/==xpc10))  xpc10 <= 13'sd2233/*2233:xpc10*/;
                  if ((13'sd2233/*2233:xpc10*/==xpc10))  xpc10 <= 13'sd2234/*2234:xpc10*/;
                  if ((13'sd2234/*2234:xpc10*/==xpc10))  xpc10 <= 13'sd2235/*2235:xpc10*/;
                  if ((13'sd2235/*2235:xpc10*/==xpc10))  xpc10 <= 13'sd1698/*1698:xpc10*/;
                  if ((13'sd2236/*2236:xpc10*/==xpc10))  xpc10 <= 13'sd2237/*2237:xpc10*/;
                  if ((13'sd2237/*2237:xpc10*/==xpc10))  xpc10 <= 13'sd2238/*2238:xpc10*/;
                  if ((13'sd2239/*2239:xpc10*/==xpc10))  xpc10 <= 13'sd2240/*2240:xpc10*/;
                  if ((13'sd2240/*2240:xpc10*/==xpc10))  xpc10 <= 13'sd2241/*2241:xpc10*/;
                  if ((13'sd2241/*2241:xpc10*/==xpc10))  xpc10 <= 13'sd2242/*2242:xpc10*/;
                  if ((13'sd2242/*2242:xpc10*/==xpc10))  xpc10 <= 13'sd2081/*2081:xpc10*/;
                  if ((13'sd2243/*2243:xpc10*/==xpc10))  xpc10 <= 13'sd2244/*2244:xpc10*/;
                  if ((13'sd2244/*2244:xpc10*/==xpc10))  xpc10 <= 13'sd2245/*2245:xpc10*/;
                  if ((13'sd2245/*2245:xpc10*/==xpc10))  xpc10 <= 13'sd2246/*2246:xpc10*/;
                  if ((13'sd2246/*2246:xpc10*/==xpc10))  xpc10 <= 13'sd2247/*2247:xpc10*/;
                  if ((13'sd2247/*2247:xpc10*/==xpc10))  xpc10 <= 13'sd2248/*2248:xpc10*/;
                  if ((13'sd2248/*2248:xpc10*/==xpc10))  xpc10 <= 13'sd2249/*2249:xpc10*/;
                  if ((13'sd2251/*2251:xpc10*/==xpc10))  xpc10 <= 13'sd1641/*1641:xpc10*/;
                  if ((13'sd2252/*2252:xpc10*/==xpc10))  xpc10 <= 13'sd2253/*2253:xpc10*/;
                  if ((13'sd2253/*2253:xpc10*/==xpc10))  xpc10 <= 13'sd2254/*2254:xpc10*/;
                  if ((13'sd2255/*2255:xpc10*/==xpc10))  xpc10 <= 13'sd798/*798:xpc10*/;
                  if ((13'sd2256/*2256:xpc10*/==xpc10))  xpc10 <= 13'sd2257/*2257:xpc10*/;
                  if ((13'sd2257/*2257:xpc10*/==xpc10))  xpc10 <= 13'sd2258/*2258:xpc10*/;
                  if ((13'sd2259/*2259:xpc10*/==xpc10))  xpc10 <= 13'sd789/*789:xpc10*/;
                  if ((13'sd2260/*2260:xpc10*/==xpc10))  xpc10 <= 13'sd2261/*2261:xpc10*/;
                  if ((13'sd2261/*2261:xpc10*/==xpc10))  xpc10 <= 13'sd2262/*2262:xpc10*/;
                  if ((13'sd2263/*2263:xpc10*/==xpc10))  xpc10 <= 13'sd2264/*2264:xpc10*/;
                  if ((13'sd2264/*2264:xpc10*/==xpc10))  xpc10 <= 13'sd2265/*2265:xpc10*/;
                  if ((13'sd2265/*2265:xpc10*/==xpc10))  xpc10 <= 13'sd2266/*2266:xpc10*/;
                  if ((13'sd2267/*2267:xpc10*/==xpc10))  xpc10 <= 13'sd776/*776:xpc10*/;
                  if ((13'sd2268/*2268:xpc10*/==xpc10))  xpc10 <= 13'sd2269/*2269:xpc10*/;
                  if ((13'sd2269/*2269:xpc10*/==xpc10))  xpc10 <= 13'sd2270/*2270:xpc10*/;
                  if ((13'sd2271/*2271:xpc10*/==xpc10))  xpc10 <= 13'sd2272/*2272:xpc10*/;
                  if ((13'sd2272/*2272:xpc10*/==xpc10))  xpc10 <= 13'sd2273/*2273:xpc10*/;
                  if ((13'sd2273/*2273:xpc10*/==xpc10))  xpc10 <= 13'sd2274/*2274:xpc10*/;
                  if ((13'sd2275/*2275:xpc10*/==xpc10))  xpc10 <= 13'sd776/*776:xpc10*/;
                  if ((13'sd2276/*2276:xpc10*/==xpc10))  xpc10 <= 13'sd2277/*2277:xpc10*/;
                  if ((13'sd2277/*2277:xpc10*/==xpc10))  xpc10 <= 13'sd2278/*2278:xpc10*/;
                  if ((13'sd2279/*2279:xpc10*/==xpc10))  xpc10 <= 13'sd776/*776:xpc10*/;
                  if ((13'sd2280/*2280:xpc10*/==xpc10))  xpc10 <= 13'sd2281/*2281:xpc10*/;
                  if ((13'sd2281/*2281:xpc10*/==xpc10))  xpc10 <= 13'sd2282/*2282:xpc10*/;
                  if ((13'sd2283/*2283:xpc10*/==xpc10))  xpc10 <= 13'sd757/*757:xpc10*/;
                  if ((13'sd2284/*2284:xpc10*/==xpc10))  xpc10 <= 13'sd2285/*2285:xpc10*/;
                  if ((13'sd2285/*2285:xpc10*/==xpc10))  xpc10 <= 13'sd2286/*2286:xpc10*/;
                  if ((13'sd2287/*2287:xpc10*/==xpc10))  xpc10 <= 13'sd747/*747:xpc10*/;
                  if ((13'sd2288/*2288:xpc10*/==xpc10))  xpc10 <= 13'sd2289/*2289:xpc10*/;
                  if ((13'sd2289/*2289:xpc10*/==xpc10))  xpc10 <= 13'sd2290/*2290:xpc10*/;
                  if ((13'sd2291/*2291:xpc10*/==xpc10))  xpc10 <= 13'sd2292/*2292:xpc10*/;
                  if ((13'sd2292/*2292:xpc10*/==xpc10))  xpc10 <= 13'sd2293/*2293:xpc10*/;
                  if ((13'sd2293/*2293:xpc10*/==xpc10))  xpc10 <= 13'sd2294/*2294:xpc10*/;
                  if ((13'sd2295/*2295:xpc10*/==xpc10))  xpc10 <= 13'sd2296/*2296:xpc10*/;
                  if ((13'sd2296/*2296:xpc10*/==xpc10))  xpc10 <= 13'sd2297/*2297:xpc10*/;
                  if ((13'sd2297/*2297:xpc10*/==xpc10))  xpc10 <= 13'sd2298/*2298:xpc10*/;
                  if ((13'sd2301/*2301:xpc10*/==xpc10))  xpc10 <= 13'sd2302/*2302:xpc10*/;
                  if ((13'sd2302/*2302:xpc10*/==xpc10))  xpc10 <= 13'sd2303/*2303:xpc10*/;
                  if ((13'sd2303/*2303:xpc10*/==xpc10))  xpc10 <= 13'sd2304/*2304:xpc10*/;
                  if ((13'sd2305/*2305:xpc10*/==xpc10))  xpc10 <= 13'sd2306/*2306:xpc10*/;
                  if ((13'sd2306/*2306:xpc10*/==xpc10))  xpc10 <= 13'sd2307/*2307:xpc10*/;
                  if ((13'sd2307/*2307:xpc10*/==xpc10))  xpc10 <= 13'sd2308/*2308:xpc10*/;
                  if ((13'sd2311/*2311:xpc10*/==xpc10))  xpc10 <= 13'sd2312/*2312:xpc10*/;
                  if ((13'sd2312/*2312:xpc10*/==xpc10))  xpc10 <= 13'sd2313/*2313:xpc10*/;
                  if ((13'sd2313/*2313:xpc10*/==xpc10))  xpc10 <= 13'sd2314/*2314:xpc10*/;
                  if ((13'sd2315/*2315:xpc10*/==xpc10))  xpc10 <= 13'sd2316/*2316:xpc10*/;
                  if ((13'sd2316/*2316:xpc10*/==xpc10))  xpc10 <= 13'sd2317/*2317:xpc10*/;
                  if ((13'sd2317/*2317:xpc10*/==xpc10))  xpc10 <= 13'sd2318/*2318:xpc10*/;
                  if ((13'sd2322/*2322:xpc10*/==xpc10))  xpc10 <= 13'sd2323/*2323:xpc10*/;
                  if ((13'sd2323/*2323:xpc10*/==xpc10))  xpc10 <= 13'sd2324/*2324:xpc10*/;
                  if ((13'sd2324/*2324:xpc10*/==xpc10))  xpc10 <= 13'sd2325/*2325:xpc10*/;
                  if ((13'sd2325/*2325:xpc10*/==xpc10))  xpc10 <= 13'sd2326/*2326:xpc10*/;
                  if ((13'sd2326/*2326:xpc10*/==xpc10))  xpc10 <= 13'sd2327/*2327:xpc10*/;
                  if ((13'sd2327/*2327:xpc10*/==xpc10))  xpc10 <= 13'sd2328/*2328:xpc10*/;
                  if ((13'sd2328/*2328:xpc10*/==xpc10))  xpc10 <= 13'sd2329/*2329:xpc10*/;
                  if ((13'sd2330/*2330:xpc10*/==xpc10))  xpc10 <= 13'sd2331/*2331:xpc10*/;
                  if ((13'sd2331/*2331:xpc10*/==xpc10))  xpc10 <= 13'sd2332/*2332:xpc10*/;
                  if ((13'sd2332/*2332:xpc10*/==xpc10))  xpc10 <= 13'sd2333/*2333:xpc10*/;
                  if ((13'sd2334/*2334:xpc10*/==xpc10))  xpc10 <= 13'sd2335/*2335:xpc10*/;
                  if ((13'sd2335/*2335:xpc10*/==xpc10))  xpc10 <= 13'sd2336/*2336:xpc10*/;
                  if ((13'sd2336/*2336:xpc10*/==xpc10))  xpc10 <= 13'sd2337/*2337:xpc10*/;
                  if ((13'sd2338/*2338:xpc10*/==xpc10))  xpc10 <= 13'sd780/*780:xpc10*/;
                  if ((13'sd2339/*2339:xpc10*/==xpc10))  xpc10 <= 13'sd2340/*2340:xpc10*/;
                  if ((13'sd2340/*2340:xpc10*/==xpc10))  xpc10 <= 13'sd2341/*2341:xpc10*/;
                  if ((13'sd2342/*2342:xpc10*/==xpc10))  xpc10 <= 13'sd2343/*2343:xpc10*/;
                  if ((13'sd2343/*2343:xpc10*/==xpc10))  xpc10 <= 13'sd2344/*2344:xpc10*/;
                  if ((13'sd2344/*2344:xpc10*/==xpc10))  xpc10 <= 13'sd2345/*2345:xpc10*/;
                  if ((13'sd2346/*2346:xpc10*/==xpc10))  xpc10 <= 13'sd2335/*2335:xpc10*/;
                  if ((13'sd2347/*2347:xpc10*/==xpc10))  xpc10 <= 13'sd2348/*2348:xpc10*/;
                  if ((13'sd2348/*2348:xpc10*/==xpc10))  xpc10 <= 13'sd2349/*2349:xpc10*/;
                  if ((13'sd2350/*2350:xpc10*/==xpc10))  xpc10 <= 13'sd2351/*2351:xpc10*/;
                  if ((13'sd2351/*2351:xpc10*/==xpc10))  xpc10 <= 13'sd2352/*2352:xpc10*/;
                  if ((13'sd2352/*2352:xpc10*/==xpc10))  xpc10 <= 13'sd2353/*2353:xpc10*/;
                  if ((13'sd2354/*2354:xpc10*/==xpc10))  xpc10 <= 13'sd2335/*2335:xpc10*/;
                  if ((13'sd2355/*2355:xpc10*/==xpc10))  xpc10 <= 13'sd2356/*2356:xpc10*/;
                  if ((13'sd2356/*2356:xpc10*/==xpc10))  xpc10 <= 13'sd2357/*2357:xpc10*/;
                  if ((13'sd2358/*2358:xpc10*/==xpc10))  xpc10 <= 13'sd2335/*2335:xpc10*/;
                  if ((13'sd2359/*2359:xpc10*/==xpc10))  xpc10 <= 13'sd2360/*2360:xpc10*/;
                  if ((13'sd2360/*2360:xpc10*/==xpc10))  xpc10 <= 13'sd2361/*2361:xpc10*/;
                  if ((13'sd2362/*2362:xpc10*/==xpc10))  xpc10 <= 13'sd2316/*2316:xpc10*/;
                  if ((13'sd2363/*2363:xpc10*/==xpc10))  xpc10 <= 13'sd2364/*2364:xpc10*/;
                  if ((13'sd2364/*2364:xpc10*/==xpc10))  xpc10 <= 13'sd2365/*2365:xpc10*/;
                  if ((13'sd2366/*2366:xpc10*/==xpc10))  xpc10 <= 13'sd2306/*2306:xpc10*/;
                  if ((13'sd2367/*2367:xpc10*/==xpc10))  xpc10 <= 13'sd2368/*2368:xpc10*/;
                  if ((13'sd2368/*2368:xpc10*/==xpc10))  xpc10 <= 13'sd2369/*2369:xpc10*/;
                  if ((13'sd2369/*2369:xpc10*/==xpc10))  xpc10 <= 13'sd2370/*2370:xpc10*/;
                  if ((13'sd2371/*2371:xpc10*/==xpc10))  xpc10 <= 13'sd780/*780:xpc10*/;
                  if ((13'sd2372/*2372:xpc10*/==xpc10))  xpc10 <= 13'sd2373/*2373:xpc10*/;
                  if ((13'sd2373/*2373:xpc10*/==xpc10))  xpc10 <= 13'sd2374/*2374:xpc10*/;
                  if ((13'sd2375/*2375:xpc10*/==xpc10))  xpc10 <= 13'sd2376/*2376:xpc10*/;
                  if ((13'sd2376/*2376:xpc10*/==xpc10))  xpc10 <= 13'sd2377/*2377:xpc10*/;
                  if ((13'sd2377/*2377:xpc10*/==xpc10))  xpc10 <= 13'sd2378/*2378:xpc10*/;
                  if ((13'sd2379/*2379:xpc10*/==xpc10))  xpc10 <= 13'sd2380/*2380:xpc10*/;
                  if ((13'sd2380/*2380:xpc10*/==xpc10))  xpc10 <= 13'sd2381/*2381:xpc10*/;
                  if ((13'sd2381/*2381:xpc10*/==xpc10))  xpc10 <= 13'sd2382/*2382:xpc10*/;
                  if ((13'sd2383/*2383:xpc10*/==xpc10))  xpc10 <= 13'sd780/*780:xpc10*/;
                  if ((13'sd2384/*2384:xpc10*/==xpc10))  xpc10 <= 13'sd2385/*2385:xpc10*/;
                  if ((13'sd2385/*2385:xpc10*/==xpc10))  xpc10 <= 13'sd2386/*2386:xpc10*/;
                  if ((13'sd2387/*2387:xpc10*/==xpc10))  xpc10 <= 13'sd2380/*2380:xpc10*/;
                  if ((13'sd2388/*2388:xpc10*/==xpc10))  xpc10 <= 13'sd2389/*2389:xpc10*/;
                  if ((13'sd2389/*2389:xpc10*/==xpc10))  xpc10 <= 13'sd2390/*2390:xpc10*/;
                  if ((13'sd2391/*2391:xpc10*/==xpc10))  xpc10 <= 13'sd2392/*2392:xpc10*/;
                  if ((13'sd2392/*2392:xpc10*/==xpc10))  xpc10 <= 13'sd2393/*2393:xpc10*/;
                  if ((13'sd2393/*2393:xpc10*/==xpc10))  xpc10 <= 13'sd2394/*2394:xpc10*/;
                  if ((13'sd2395/*2395:xpc10*/==xpc10))  xpc10 <= 13'sd2396/*2396:xpc10*/;
                  if ((13'sd2396/*2396:xpc10*/==xpc10))  xpc10 <= 13'sd2397/*2397:xpc10*/;
                  if ((13'sd2397/*2397:xpc10*/==xpc10))  xpc10 <= 13'sd2398/*2398:xpc10*/;
                  if ((13'sd2401/*2401:xpc10*/==xpc10))  xpc10 <= 13'sd2402/*2402:xpc10*/;
                  if ((13'sd2402/*2402:xpc10*/==xpc10))  xpc10 <= 13'sd2403/*2403:xpc10*/;
                  if ((13'sd2403/*2403:xpc10*/==xpc10))  xpc10 <= 13'sd2404/*2404:xpc10*/;
                  if ((13'sd2405/*2405:xpc10*/==xpc10))  xpc10 <= 13'sd2406/*2406:xpc10*/;
                  if ((13'sd2406/*2406:xpc10*/==xpc10))  xpc10 <= 13'sd2407/*2407:xpc10*/;
                  if ((13'sd2407/*2407:xpc10*/==xpc10))  xpc10 <= 13'sd2408/*2408:xpc10*/;
                  if ((13'sd2411/*2411:xpc10*/==xpc10))  xpc10 <= 13'sd2412/*2412:xpc10*/;
                  if ((13'sd2412/*2412:xpc10*/==xpc10))  xpc10 <= 13'sd2413/*2413:xpc10*/;
                  if ((13'sd2413/*2413:xpc10*/==xpc10))  xpc10 <= 13'sd2414/*2414:xpc10*/;
                  if ((13'sd2415/*2415:xpc10*/==xpc10))  xpc10 <= 13'sd2416/*2416:xpc10*/;
                  if ((13'sd2416/*2416:xpc10*/==xpc10))  xpc10 <= 13'sd2417/*2417:xpc10*/;
                  if ((13'sd2417/*2417:xpc10*/==xpc10))  xpc10 <= 13'sd2418/*2418:xpc10*/;
                  if ((13'sd2422/*2422:xpc10*/==xpc10))  xpc10 <= 13'sd2423/*2423:xpc10*/;
                  if ((13'sd2423/*2423:xpc10*/==xpc10))  xpc10 <= 13'sd2424/*2424:xpc10*/;
                  if ((13'sd2424/*2424:xpc10*/==xpc10))  xpc10 <= 13'sd2425/*2425:xpc10*/;
                  if ((13'sd2425/*2425:xpc10*/==xpc10))  xpc10 <= 13'sd2426/*2426:xpc10*/;
                  if ((13'sd2426/*2426:xpc10*/==xpc10))  xpc10 <= 13'sd2427/*2427:xpc10*/;
                  if ((13'sd2427/*2427:xpc10*/==xpc10))  xpc10 <= 13'sd2428/*2428:xpc10*/;
                  if ((13'sd2428/*2428:xpc10*/==xpc10))  xpc10 <= 13'sd2429/*2429:xpc10*/;
                  if ((13'sd2430/*2430:xpc10*/==xpc10))  xpc10 <= 13'sd2431/*2431:xpc10*/;
                  if ((13'sd2431/*2431:xpc10*/==xpc10))  xpc10 <= 13'sd2432/*2432:xpc10*/;
                  if ((13'sd2432/*2432:xpc10*/==xpc10))  xpc10 <= 13'sd2433/*2433:xpc10*/;
                  if ((13'sd2434/*2434:xpc10*/==xpc10))  xpc10 <= 13'sd2435/*2435:xpc10*/;
                  if ((13'sd2435/*2435:xpc10*/==xpc10))  xpc10 <= 13'sd2436/*2436:xpc10*/;
                  if ((13'sd2436/*2436:xpc10*/==xpc10))  xpc10 <= 13'sd2437/*2437:xpc10*/;
                  if ((13'sd2438/*2438:xpc10*/==xpc10))  xpc10 <= 13'sd780/*780:xpc10*/;
                  if ((13'sd2439/*2439:xpc10*/==xpc10))  xpc10 <= 13'sd2440/*2440:xpc10*/;
                  if ((13'sd2440/*2440:xpc10*/==xpc10))  xpc10 <= 13'sd2441/*2441:xpc10*/;
                  if ((13'sd2442/*2442:xpc10*/==xpc10))  xpc10 <= 13'sd2443/*2443:xpc10*/;
                  if ((13'sd2443/*2443:xpc10*/==xpc10))  xpc10 <= 13'sd2444/*2444:xpc10*/;
                  if ((13'sd2444/*2444:xpc10*/==xpc10))  xpc10 <= 13'sd2445/*2445:xpc10*/;
                  if ((13'sd2446/*2446:xpc10*/==xpc10))  xpc10 <= 13'sd2435/*2435:xpc10*/;
                  if ((13'sd2447/*2447:xpc10*/==xpc10))  xpc10 <= 13'sd2448/*2448:xpc10*/;
                  if ((13'sd2448/*2448:xpc10*/==xpc10))  xpc10 <= 13'sd2449/*2449:xpc10*/;
                  if ((13'sd2450/*2450:xpc10*/==xpc10))  xpc10 <= 13'sd2451/*2451:xpc10*/;
                  if ((13'sd2451/*2451:xpc10*/==xpc10))  xpc10 <= 13'sd2452/*2452:xpc10*/;
                  if ((13'sd2452/*2452:xpc10*/==xpc10))  xpc10 <= 13'sd2453/*2453:xpc10*/;
                  if ((13'sd2454/*2454:xpc10*/==xpc10))  xpc10 <= 13'sd2435/*2435:xpc10*/;
                  if ((13'sd2455/*2455:xpc10*/==xpc10))  xpc10 <= 13'sd2456/*2456:xpc10*/;
                  if ((13'sd2456/*2456:xpc10*/==xpc10))  xpc10 <= 13'sd2457/*2457:xpc10*/;
                  if ((13'sd2458/*2458:xpc10*/==xpc10))  xpc10 <= 13'sd2435/*2435:xpc10*/;
                  if ((13'sd2459/*2459:xpc10*/==xpc10))  xpc10 <= 13'sd2460/*2460:xpc10*/;
                  if ((13'sd2460/*2460:xpc10*/==xpc10))  xpc10 <= 13'sd2461/*2461:xpc10*/;
                  if ((13'sd2462/*2462:xpc10*/==xpc10))  xpc10 <= 13'sd2416/*2416:xpc10*/;
                  if ((13'sd2463/*2463:xpc10*/==xpc10))  xpc10 <= 13'sd2464/*2464:xpc10*/;
                  if ((13'sd2464/*2464:xpc10*/==xpc10))  xpc10 <= 13'sd2465/*2465:xpc10*/;
                  if ((13'sd2466/*2466:xpc10*/==xpc10))  xpc10 <= 13'sd2406/*2406:xpc10*/;
                  if ((13'sd2467/*2467:xpc10*/==xpc10))  xpc10 <= 13'sd2468/*2468:xpc10*/;
                  if ((13'sd2468/*2468:xpc10*/==xpc10))  xpc10 <= 13'sd2469/*2469:xpc10*/;
                  if ((13'sd2470/*2470:xpc10*/==xpc10))  xpc10 <= 13'sd2471/*2471:xpc10*/;
                  if ((13'sd2471/*2471:xpc10*/==xpc10))  xpc10 <= 13'sd2472/*2472:xpc10*/;
                  if ((13'sd2472/*2472:xpc10*/==xpc10))  xpc10 <= 13'sd2473/*2473:xpc10*/;
                  if ((13'sd2474/*2474:xpc10*/==xpc10))  xpc10 <= 13'sd2475/*2475:xpc10*/;
                  if ((13'sd2475/*2475:xpc10*/==xpc10))  xpc10 <= 13'sd2476/*2476:xpc10*/;
                  if ((13'sd2476/*2476:xpc10*/==xpc10))  xpc10 <= 13'sd2477/*2477:xpc10*/;
                  if ((13'sd2478/*2478:xpc10*/==xpc10))  xpc10 <= 13'sd780/*780:xpc10*/;
                  if ((13'sd2479/*2479:xpc10*/==xpc10))  xpc10 <= 13'sd2480/*2480:xpc10*/;
                  if ((13'sd2480/*2480:xpc10*/==xpc10))  xpc10 <= 13'sd2481/*2481:xpc10*/;
                  if ((13'sd2482/*2482:xpc10*/==xpc10))  xpc10 <= 13'sd2475/*2475:xpc10*/;
                  if ((13'sd2483/*2483:xpc10*/==xpc10))  xpc10 <= 13'sd2484/*2484:xpc10*/;
                  if ((13'sd2484/*2484:xpc10*/==xpc10))  xpc10 <= 13'sd2485/*2485:xpc10*/;
                  if ((13'sd2486/*2486:xpc10*/==xpc10))  xpc10 <= 13'sd2487/*2487:xpc10*/;
                  if ((13'sd2487/*2487:xpc10*/==xpc10))  xpc10 <= 13'sd2488/*2488:xpc10*/;
                  if ((13'sd2488/*2488:xpc10*/==xpc10))  xpc10 <= 13'sd2489/*2489:xpc10*/;
                  if ((13'sd2490/*2490:xpc10*/==xpc10))  xpc10 <= 13'sd2491/*2491:xpc10*/;
                  if ((13'sd2491/*2491:xpc10*/==xpc10))  xpc10 <= 13'sd2492/*2492:xpc10*/;
                  if ((13'sd2492/*2492:xpc10*/==xpc10))  xpc10 <= 13'sd2493/*2493:xpc10*/;
                  if ((13'sd2494/*2494:xpc10*/==xpc10))  xpc10 <= 13'sd2495/*2495:xpc10*/;
                  if ((13'sd2495/*2495:xpc10*/==xpc10))  xpc10 <= 13'sd2496/*2496:xpc10*/;
                  if ((13'sd2496/*2496:xpc10*/==xpc10))  xpc10 <= 13'sd2497/*2497:xpc10*/;
                  if ((13'sd2498/*2498:xpc10*/==xpc10))  xpc10 <= 13'sd2499/*2499:xpc10*/;
                  if ((13'sd2499/*2499:xpc10*/==xpc10))  xpc10 <= 13'sd2500/*2500:xpc10*/;
                  if ((13'sd2500/*2500:xpc10*/==xpc10))  xpc10 <= 13'sd2501/*2501:xpc10*/;
                  if ((13'sd2501/*2501:xpc10*/==xpc10))  xpc10 <= 13'sd2502/*2502:xpc10*/;
                  if ((13'sd2503/*2503:xpc10*/==xpc10))  xpc10 <= 13'sd780/*780:xpc10*/;
                  if ((13'sd2504/*2504:xpc10*/==xpc10))  xpc10 <= 13'sd2505/*2505:xpc10*/;
                  if ((13'sd2505/*2505:xpc10*/==xpc10))  xpc10 <= 13'sd2506/*2506:xpc10*/;
                  if ((13'sd2506/*2506:xpc10*/==xpc10))  xpc10 <= 13'sd2507/*2507:xpc10*/;
                  if ((13'sd2508/*2508:xpc10*/==xpc10))  xpc10 <= 13'sd2509/*2509:xpc10*/;
                  if ((13'sd2509/*2509:xpc10*/==xpc10))  xpc10 <= 13'sd2510/*2510:xpc10*/;
                  if ((13'sd2510/*2510:xpc10*/==xpc10))  xpc10 <= 13'sd2511/*2511:xpc10*/;
                  if ((13'sd2512/*2512:xpc10*/==xpc10))  xpc10 <= 13'sd2513/*2513:xpc10*/;
                  if ((13'sd2513/*2513:xpc10*/==xpc10))  xpc10 <= 13'sd2514/*2514:xpc10*/;
                  if ((13'sd2514/*2514:xpc10*/==xpc10))  xpc10 <= 13'sd2515/*2515:xpc10*/;
                  if ((13'sd2516/*2516:xpc10*/==xpc10))  xpc10 <= 13'sd780/*780:xpc10*/;
                  if ((13'sd2517/*2517:xpc10*/==xpc10))  xpc10 <= 13'sd2518/*2518:xpc10*/;
                  if ((13'sd2518/*2518:xpc10*/==xpc10))  xpc10 <= 13'sd2519/*2519:xpc10*/;
                  if ((13'sd2520/*2520:xpc10*/==xpc10))  xpc10 <= 13'sd2513/*2513:xpc10*/;
                  if ((13'sd2521/*2521:xpc10*/==xpc10))  xpc10 <= 13'sd2522/*2522:xpc10*/;
                  if ((13'sd2522/*2522:xpc10*/==xpc10))  xpc10 <= 13'sd2523/*2523:xpc10*/;
                  if ((13'sd2526/*2526:xpc10*/==xpc10))  xpc10 <= 13'sd2527/*2527:xpc10*/;
                  if ((13'sd2527/*2527:xpc10*/==xpc10))  xpc10 <= 13'sd2528/*2528:xpc10*/;
                  if ((13'sd2528/*2528:xpc10*/==xpc10))  xpc10 <= 13'sd2529/*2529:xpc10*/;
                  if ((13'sd2530/*2530:xpc10*/==xpc10))  xpc10 <= 13'sd2531/*2531:xpc10*/;
                  if ((13'sd2531/*2531:xpc10*/==xpc10))  xpc10 <= 13'sd2532/*2532:xpc10*/;
                  if ((13'sd2532/*2532:xpc10*/==xpc10))  xpc10 <= 13'sd2533/*2533:xpc10*/;
                  if ((13'sd2536/*2536:xpc10*/==xpc10))  xpc10 <= 13'sd2537/*2537:xpc10*/;
                  if ((13'sd2537/*2537:xpc10*/==xpc10))  xpc10 <= 13'sd2538/*2538:xpc10*/;
                  if ((13'sd2538/*2538:xpc10*/==xpc10))  xpc10 <= 13'sd2539/*2539:xpc10*/;
                  if ((13'sd2541/*2541:xpc10*/==xpc10))  xpc10 <= 13'sd2542/*2542:xpc10*/;
                  if ((13'sd2542/*2542:xpc10*/==xpc10))  xpc10 <= 13'sd2543/*2543:xpc10*/;
                  if ((13'sd2543/*2543:xpc10*/==xpc10))  xpc10 <= 13'sd2544/*2544:xpc10*/;
                  if ((13'sd2545/*2545:xpc10*/==xpc10))  xpc10 <= 13'sd2546/*2546:xpc10*/;
                  if ((13'sd2546/*2546:xpc10*/==xpc10))  xpc10 <= 13'sd2547/*2547:xpc10*/;
                  if ((13'sd2547/*2547:xpc10*/==xpc10))  xpc10 <= 13'sd2548/*2548:xpc10*/;
                  if ((13'sd2550/*2550:xpc10*/==xpc10))  xpc10 <= 13'sd2551/*2551:xpc10*/;
                  if ((13'sd2551/*2551:xpc10*/==xpc10))  xpc10 <= 13'sd2552/*2552:xpc10*/;
                  if ((13'sd2552/*2552:xpc10*/==xpc10))  xpc10 <= 13'sd2553/*2553:xpc10*/;
                  if ((13'sd2558/*2558:xpc10*/==xpc10))  xpc10 <= 13'sd2559/*2559:xpc10*/;
                  if ((13'sd2559/*2559:xpc10*/==xpc10))  xpc10 <= 13'sd2560/*2560:xpc10*/;
                  if ((13'sd2560/*2560:xpc10*/==xpc10))  xpc10 <= 13'sd2561/*2561:xpc10*/;
                  if ((13'sd2562/*2562:xpc10*/==xpc10))  xpc10 <= 13'sd2563/*2563:xpc10*/;
                  if ((13'sd2563/*2563:xpc10*/==xpc10))  xpc10 <= 13'sd2564/*2564:xpc10*/;
                  if ((13'sd2564/*2564:xpc10*/==xpc10))  xpc10 <= 13'sd2565/*2565:xpc10*/;
                  if ((13'sd2566/*2566:xpc10*/==xpc10))  xpc10 <= 13'sd2567/*2567:xpc10*/;
                  if ((13'sd2567/*2567:xpc10*/==xpc10))  xpc10 <= 13'sd2568/*2568:xpc10*/;
                  if ((13'sd2568/*2568:xpc10*/==xpc10))  xpc10 <= 13'sd2569/*2569:xpc10*/;
                  if ((13'sd2570/*2570:xpc10*/==xpc10))  xpc10 <= 13'sd2571/*2571:xpc10*/;
                  if ((13'sd2571/*2571:xpc10*/==xpc10))  xpc10 <= 13'sd2572/*2572:xpc10*/;
                  if ((13'sd2572/*2572:xpc10*/==xpc10))  xpc10 <= 13'sd2573/*2573:xpc10*/;
                  if ((13'sd2574/*2574:xpc10*/==xpc10))  xpc10 <= 13'sd2575/*2575:xpc10*/;
                  if ((13'sd2575/*2575:xpc10*/==xpc10))  xpc10 <= 13'sd2576/*2576:xpc10*/;
                  if ((13'sd2576/*2576:xpc10*/==xpc10))  xpc10 <= 13'sd2577/*2577:xpc10*/;
                  if ((13'sd2578/*2578:xpc10*/==xpc10))  xpc10 <= 13'sd780/*780:xpc10*/;
                  if ((13'sd2579/*2579:xpc10*/==xpc10))  xpc10 <= 13'sd2580/*2580:xpc10*/;
                  if ((13'sd2580/*2580:xpc10*/==xpc10))  xpc10 <= 13'sd2581/*2581:xpc10*/;
                  if ((13'sd2582/*2582:xpc10*/==xpc10))  xpc10 <= 13'sd2575/*2575:xpc10*/;
                  if ((13'sd2583/*2583:xpc10*/==xpc10))  xpc10 <= 13'sd2584/*2584:xpc10*/;
                  if ((13'sd2584/*2584:xpc10*/==xpc10))  xpc10 <= 13'sd2585/*2585:xpc10*/;
                  if ((13'sd2588/*2588:xpc10*/==xpc10))  xpc10 <= 13'sd2589/*2589:xpc10*/;
                  if ((13'sd2589/*2589:xpc10*/==xpc10))  xpc10 <= 13'sd2590/*2590:xpc10*/;
                  if ((13'sd2590/*2590:xpc10*/==xpc10))  xpc10 <= 13'sd2591/*2591:xpc10*/;
                  if ((13'sd2592/*2592:xpc10*/==xpc10))  xpc10 <= 13'sd2593/*2593:xpc10*/;
                  if ((13'sd2593/*2593:xpc10*/==xpc10))  xpc10 <= 13'sd2594/*2594:xpc10*/;
                  if ((13'sd2594/*2594:xpc10*/==xpc10))  xpc10 <= 13'sd2595/*2595:xpc10*/;
                  if ((13'sd2598/*2598:xpc10*/==xpc10))  xpc10 <= 13'sd2599/*2599:xpc10*/;
                  if ((13'sd2599/*2599:xpc10*/==xpc10))  xpc10 <= 13'sd2600/*2600:xpc10*/;
                  if ((13'sd2600/*2600:xpc10*/==xpc10))  xpc10 <= 13'sd2601/*2601:xpc10*/;
                  if ((13'sd2603/*2603:xpc10*/==xpc10))  xpc10 <= 13'sd2604/*2604:xpc10*/;
                  if ((13'sd2604/*2604:xpc10*/==xpc10))  xpc10 <= 13'sd2605/*2605:xpc10*/;
                  if ((13'sd2605/*2605:xpc10*/==xpc10))  xpc10 <= 13'sd2606/*2606:xpc10*/;
                  if ((13'sd2607/*2607:xpc10*/==xpc10))  xpc10 <= 13'sd2608/*2608:xpc10*/;
                  if ((13'sd2608/*2608:xpc10*/==xpc10))  xpc10 <= 13'sd2609/*2609:xpc10*/;
                  if ((13'sd2609/*2609:xpc10*/==xpc10))  xpc10 <= 13'sd2610/*2610:xpc10*/;
                  if ((13'sd2612/*2612:xpc10*/==xpc10))  xpc10 <= 13'sd2613/*2613:xpc10*/;
                  if ((13'sd2613/*2613:xpc10*/==xpc10))  xpc10 <= 13'sd2614/*2614:xpc10*/;
                  if ((13'sd2614/*2614:xpc10*/==xpc10))  xpc10 <= 13'sd2615/*2615:xpc10*/;
                  if ((13'sd2620/*2620:xpc10*/==xpc10))  xpc10 <= 13'sd2621/*2621:xpc10*/;
                  if ((13'sd2621/*2621:xpc10*/==xpc10))  xpc10 <= 13'sd2622/*2622:xpc10*/;
                  if ((13'sd2622/*2622:xpc10*/==xpc10))  xpc10 <= 13'sd2623/*2623:xpc10*/;
                  if ((13'sd2627/*2627:xpc10*/==xpc10))  xpc10 <= 13'sd2628/*2628:xpc10*/;
                  if ((13'sd2628/*2628:xpc10*/==xpc10))  xpc10 <= 13'sd2629/*2629:xpc10*/;
                  if ((13'sd2629/*2629:xpc10*/==xpc10))  xpc10 <= 13'sd2630/*2630:xpc10*/;
                  if ((13'sd2632/*2632:xpc10*/==xpc10))  xpc10 <= 13'sd2633/*2633:xpc10*/;
                  if ((13'sd2633/*2633:xpc10*/==xpc10))  xpc10 <= 13'sd2634/*2634:xpc10*/;
                  if ((13'sd2634/*2634:xpc10*/==xpc10))  xpc10 <= 13'sd2635/*2635:xpc10*/;
                  if ((13'sd2636/*2636:xpc10*/==xpc10))  xpc10 <= 13'sd2637/*2637:xpc10*/;
                  if ((13'sd2637/*2637:xpc10*/==xpc10))  xpc10 <= 13'sd2638/*2638:xpc10*/;
                  if ((13'sd2638/*2638:xpc10*/==xpc10))  xpc10 <= 13'sd2639/*2639:xpc10*/;
                  if ((13'sd2640/*2640:xpc10*/==xpc10))  xpc10 <= 13'sd2641/*2641:xpc10*/;
                  if ((13'sd2641/*2641:xpc10*/==xpc10))  xpc10 <= 13'sd2642/*2642:xpc10*/;
                  if ((13'sd2642/*2642:xpc10*/==xpc10))  xpc10 <= 13'sd2643/*2643:xpc10*/;
                  if ((13'sd2645/*2645:xpc10*/==xpc10))  xpc10 <= 13'sd2646/*2646:xpc10*/;
                  if ((13'sd2646/*2646:xpc10*/==xpc10))  xpc10 <= 13'sd2647/*2647:xpc10*/;
                  if ((13'sd2647/*2647:xpc10*/==xpc10))  xpc10 <= 13'sd2648/*2648:xpc10*/;
                  if ((13'sd2658/*2658:xpc10*/==xpc10))  xpc10 <= 13'sd2659/*2659:xpc10*/;
                  if ((13'sd2659/*2659:xpc10*/==xpc10))  xpc10 <= 13'sd2660/*2660:xpc10*/;
                  if ((13'sd2660/*2660:xpc10*/==xpc10))  xpc10 <= 13'sd2661/*2661:xpc10*/;
                  if ((13'sd2661/*2661:xpc10*/==xpc10))  xpc10 <= 13'sd2662/*2662:xpc10*/;
                  if ((13'sd2662/*2662:xpc10*/==xpc10))  xpc10 <= 13'sd2663/*2663:xpc10*/;
                  if ((13'sd2663/*2663:xpc10*/==xpc10))  xpc10 <= 13'sd2664/*2664:xpc10*/;
                  if ((13'sd2664/*2664:xpc10*/==xpc10))  xpc10 <= 13'sd2665/*2665:xpc10*/;
                  if ((13'sd2665/*2665:xpc10*/==xpc10))  xpc10 <= 13'sd2666/*2666:xpc10*/;
                  if ((13'sd2670/*2670:xpc10*/==xpc10))  xpc10 <= 13'sd2671/*2671:xpc10*/;
                  if ((13'sd2671/*2671:xpc10*/==xpc10))  xpc10 <= 13'sd2672/*2672:xpc10*/;
                  if ((13'sd2672/*2672:xpc10*/==xpc10))  xpc10 <= 13'sd2673/*2673:xpc10*/;
                  if ((13'sd2675/*2675:xpc10*/==xpc10))  xpc10 <= 13'sd2676/*2676:xpc10*/;
                  if ((13'sd2676/*2676:xpc10*/==xpc10))  xpc10 <= 13'sd2677/*2677:xpc10*/;
                  if ((13'sd2677/*2677:xpc10*/==xpc10))  xpc10 <= 13'sd2678/*2678:xpc10*/;
                  if ((13'sd2685/*2685:xpc10*/==xpc10))  xpc10 <= 13'sd2686/*2686:xpc10*/;
                  if ((13'sd2686/*2686:xpc10*/==xpc10))  xpc10 <= 13'sd2687/*2687:xpc10*/;
                  if ((13'sd2687/*2687:xpc10*/==xpc10))  xpc10 <= 13'sd2688/*2688:xpc10*/;
                  if ((13'sd2690/*2690:xpc10*/==xpc10))  xpc10 <= 13'sd2691/*2691:xpc10*/;
                  if ((13'sd2691/*2691:xpc10*/==xpc10))  xpc10 <= 13'sd2692/*2692:xpc10*/;
                  if ((13'sd2692/*2692:xpc10*/==xpc10))  xpc10 <= 13'sd2693/*2693:xpc10*/;
                  if ((13'sd2701/*2701:xpc10*/==xpc10))  xpc10 <= 13'sd2702/*2702:xpc10*/;
                  if ((13'sd2702/*2702:xpc10*/==xpc10))  xpc10 <= 13'sd2703/*2703:xpc10*/;
                  if ((13'sd2703/*2703:xpc10*/==xpc10))  xpc10 <= 13'sd2704/*2704:xpc10*/;
                  if ((13'sd2706/*2706:xpc10*/==xpc10))  xpc10 <= 13'sd2707/*2707:xpc10*/;
                  if ((13'sd2707/*2707:xpc10*/==xpc10))  xpc10 <= 13'sd2708/*2708:xpc10*/;
                  if ((13'sd2708/*2708:xpc10*/==xpc10))  xpc10 <= 13'sd2709/*2709:xpc10*/;
                  if ((13'sd2710/*2710:xpc10*/==xpc10))  xpc10 <= 13'sd2711/*2711:xpc10*/;
                  if ((13'sd2711/*2711:xpc10*/==xpc10))  xpc10 <= 13'sd2712/*2712:xpc10*/;
                  if ((13'sd2712/*2712:xpc10*/==xpc10))  xpc10 <= 13'sd2713/*2713:xpc10*/;
                  if ((13'sd2714/*2714:xpc10*/==xpc10))  xpc10 <= 13'sd2715/*2715:xpc10*/;
                  if ((13'sd2715/*2715:xpc10*/==xpc10))  xpc10 <= 13'sd2716/*2716:xpc10*/;
                  if ((13'sd2716/*2716:xpc10*/==xpc10))  xpc10 <= 13'sd2717/*2717:xpc10*/;
                  if ((13'sd2721/*2721:xpc10*/==xpc10))  xpc10 <= 13'sd2722/*2722:xpc10*/;
                  if ((13'sd2722/*2722:xpc10*/==xpc10))  xpc10 <= 13'sd2723/*2723:xpc10*/;
                  if ((13'sd2723/*2723:xpc10*/==xpc10))  xpc10 <= 13'sd2724/*2724:xpc10*/;
                  if ((13'sd2726/*2726:xpc10*/==xpc10))  xpc10 <= 13'sd2727/*2727:xpc10*/;
                  if ((13'sd2727/*2727:xpc10*/==xpc10))  xpc10 <= 13'sd2728/*2728:xpc10*/;
                  if ((13'sd2728/*2728:xpc10*/==xpc10))  xpc10 <= 13'sd2729/*2729:xpc10*/;
                  if ((13'sd2730/*2730:xpc10*/==xpc10))  xpc10 <= 13'sd2731/*2731:xpc10*/;
                  if ((13'sd2731/*2731:xpc10*/==xpc10))  xpc10 <= 13'sd2732/*2732:xpc10*/;
                  if ((13'sd2732/*2732:xpc10*/==xpc10))  xpc10 <= 13'sd2733/*2733:xpc10*/;
                  if ((13'sd2735/*2735:xpc10*/==xpc10))  xpc10 <= 13'sd2736/*2736:xpc10*/;
                  if ((13'sd2736/*2736:xpc10*/==xpc10))  xpc10 <= 13'sd2737/*2737:xpc10*/;
                  if ((13'sd2738/*2738:xpc10*/==xpc10))  xpc10 <= 13'sd2739/*2739:xpc10*/;
                  if ((13'sd2739/*2739:xpc10*/==xpc10))  xpc10 <= 13'sd2740/*2740:xpc10*/;
                  if ((13'sd2740/*2740:xpc10*/==xpc10))  xpc10 <= 13'sd2741/*2741:xpc10*/;
                  if ((13'sd2743/*2743:xpc10*/==xpc10))  xpc10 <= 13'sd2744/*2744:xpc10*/;
                  if ((13'sd2744/*2744:xpc10*/==xpc10))  xpc10 <= 13'sd2745/*2745:xpc10*/;
                  if ((13'sd2745/*2745:xpc10*/==xpc10))  xpc10 <= 13'sd2746/*2746:xpc10*/;
                  if ((13'sd2747/*2747:xpc10*/==xpc10))  xpc10 <= 13'sd2748/*2748:xpc10*/;
                  if ((13'sd2748/*2748:xpc10*/==xpc10))  xpc10 <= 13'sd2749/*2749:xpc10*/;
                  if ((13'sd2749/*2749:xpc10*/==xpc10))  xpc10 <= 13'sd2750/*2750:xpc10*/;
                  if ((13'sd2751/*2751:xpc10*/==xpc10))  xpc10 <= 13'sd2752/*2752:xpc10*/;
                  if ((13'sd2752/*2752:xpc10*/==xpc10))  xpc10 <= 13'sd2753/*2753:xpc10*/;
                  if ((13'sd2753/*2753:xpc10*/==xpc10))  xpc10 <= 13'sd2754/*2754:xpc10*/;
                  if ((13'sd2755/*2755:xpc10*/==xpc10))  xpc10 <= 13'sd2756/*2756:xpc10*/;
                  if ((13'sd2756/*2756:xpc10*/==xpc10))  xpc10 <= 13'sd2757/*2757:xpc10*/;
                  if ((13'sd2757/*2757:xpc10*/==xpc10))  xpc10 <= 13'sd2758/*2758:xpc10*/;
                  if ((13'sd2758/*2758:xpc10*/==xpc10))  xpc10 <= 13'sd2759/*2759:xpc10*/;
                  if ((13'sd2760/*2760:xpc10*/==xpc10))  xpc10 <= 13'sd2761/*2761:xpc10*/;
                  if ((13'sd2761/*2761:xpc10*/==xpc10))  xpc10 <= 13'sd2762/*2762:xpc10*/;
                  if ((13'sd2762/*2762:xpc10*/==xpc10))  xpc10 <= 13'sd2763/*2763:xpc10*/;
                  if ((13'sd2764/*2764:xpc10*/==xpc10))  xpc10 <= 13'sd2765/*2765:xpc10*/;
                  if ((13'sd2765/*2765:xpc10*/==xpc10))  xpc10 <= 13'sd2766/*2766:xpc10*/;
                  if ((13'sd2766/*2766:xpc10*/==xpc10))  xpc10 <= 13'sd2767/*2767:xpc10*/;
                  if ((13'sd2771/*2771:xpc10*/==xpc10))  xpc10 <= 13'sd2772/*2772:xpc10*/;
                  if ((13'sd2772/*2772:xpc10*/==xpc10))  xpc10 <= 13'sd2773/*2773:xpc10*/;
                  if ((13'sd2773/*2773:xpc10*/==xpc10))  xpc10 <= 13'sd2774/*2774:xpc10*/;
                  if ((13'sd2776/*2776:xpc10*/==xpc10))  xpc10 <= 13'sd2777/*2777:xpc10*/;
                  if ((13'sd2777/*2777:xpc10*/==xpc10))  xpc10 <= 13'sd2778/*2778:xpc10*/;
                  if ((13'sd2778/*2778:xpc10*/==xpc10))  xpc10 <= 13'sd2779/*2779:xpc10*/;
                  if ((13'sd2780/*2780:xpc10*/==xpc10))  xpc10 <= 13'sd2781/*2781:xpc10*/;
                  if ((13'sd2781/*2781:xpc10*/==xpc10))  xpc10 <= 13'sd2782/*2782:xpc10*/;
                  if ((13'sd2782/*2782:xpc10*/==xpc10))  xpc10 <= 13'sd2783/*2783:xpc10*/;
                  if ((13'sd2784/*2784:xpc10*/==xpc10))  xpc10 <= 13'sd780/*780:xpc10*/;
                  if ((13'sd2785/*2785:xpc10*/==xpc10))  xpc10 <= 13'sd2786/*2786:xpc10*/;
                  if ((13'sd2786/*2786:xpc10*/==xpc10))  xpc10 <= 13'sd2787/*2787:xpc10*/;
                  if ((13'sd2789/*2789:xpc10*/==xpc10))  xpc10 <= 13'sd2777/*2777:xpc10*/;
                  if ((13'sd2790/*2790:xpc10*/==xpc10))  xpc10 <= 13'sd2791/*2791:xpc10*/;
                  if ((13'sd2791/*2791:xpc10*/==xpc10))  xpc10 <= 13'sd2792/*2792:xpc10*/;
                  if ((13'sd2793/*2793:xpc10*/==xpc10))  xpc10 <= 13'sd2765/*2765:xpc10*/;
                  if ((13'sd2794/*2794:xpc10*/==xpc10))  xpc10 <= 13'sd2795/*2795:xpc10*/;
                  if ((13'sd2795/*2795:xpc10*/==xpc10))  xpc10 <= 13'sd2796/*2796:xpc10*/;
                  if ((13'sd2797/*2797:xpc10*/==xpc10))  xpc10 <= 13'sd2798/*2798:xpc10*/;
                  if ((13'sd2798/*2798:xpc10*/==xpc10))  xpc10 <= 13'sd2799/*2799:xpc10*/;
                  if ((13'sd2799/*2799:xpc10*/==xpc10))  xpc10 <= 13'sd2800/*2800:xpc10*/;
                  if ((13'sd2800/*2800:xpc10*/==xpc10))  xpc10 <= 13'sd2801/*2801:xpc10*/;
                  if ((13'sd2802/*2802:xpc10*/==xpc10))  xpc10 <= 13'sd2803/*2803:xpc10*/;
                  if ((13'sd2803/*2803:xpc10*/==xpc10))  xpc10 <= 13'sd2804/*2804:xpc10*/;
                  if ((13'sd2804/*2804:xpc10*/==xpc10))  xpc10 <= 13'sd2805/*2805:xpc10*/;
                  if ((13'sd2806/*2806:xpc10*/==xpc10))  xpc10 <= 13'sd2807/*2807:xpc10*/;
                  if ((13'sd2807/*2807:xpc10*/==xpc10))  xpc10 <= 13'sd2808/*2808:xpc10*/;
                  if ((13'sd2808/*2808:xpc10*/==xpc10))  xpc10 <= 13'sd2809/*2809:xpc10*/;
                  if ((13'sd2812/*2812:xpc10*/==xpc10))  xpc10 <= 13'sd2813/*2813:xpc10*/;
                  if ((13'sd2813/*2813:xpc10*/==xpc10))  xpc10 <= 13'sd2814/*2814:xpc10*/;
                  if ((13'sd2814/*2814:xpc10*/==xpc10))  xpc10 <= 13'sd2815/*2815:xpc10*/;
                  if ((13'sd2816/*2816:xpc10*/==xpc10))  xpc10 <= 13'sd2817/*2817:xpc10*/;
                  if ((13'sd2817/*2817:xpc10*/==xpc10))  xpc10 <= 13'sd2818/*2818:xpc10*/;
                  if ((13'sd2818/*2818:xpc10*/==xpc10))  xpc10 <= 13'sd2819/*2819:xpc10*/;
                  if ((13'sd2819/*2819:xpc10*/==xpc10))  xpc10 <= 13'sd2820/*2820:xpc10*/;
                  if ((13'sd2820/*2820:xpc10*/==xpc10))  xpc10 <= 13'sd2821/*2821:xpc10*/;
                  if ((13'sd2821/*2821:xpc10*/==xpc10))  xpc10 <= 13'sd2822/*2822:xpc10*/;
                  if ((13'sd2822/*2822:xpc10*/==xpc10))  xpc10 <= 13'sd2823/*2823:xpc10*/;
                  if ((13'sd2824/*2824:xpc10*/==xpc10))  xpc10 <= 13'sd2825/*2825:xpc10*/;
                  if ((13'sd2825/*2825:xpc10*/==xpc10))  xpc10 <= 13'sd2826/*2826:xpc10*/;
                  if ((13'sd2826/*2826:xpc10*/==xpc10))  xpc10 <= 13'sd2827/*2827:xpc10*/;
                  if ((13'sd2827/*2827:xpc10*/==xpc10))  xpc10 <= 13'sd2828/*2828:xpc10*/;
                  if ((13'sd2828/*2828:xpc10*/==xpc10))  xpc10 <= 13'sd2829/*2829:xpc10*/;
                  if ((13'sd2829/*2829:xpc10*/==xpc10))  xpc10 <= 13'sd2830/*2830:xpc10*/;
                  if ((13'sd2830/*2830:xpc10*/==xpc10))  xpc10 <= 13'sd2831/*2831:xpc10*/;
                  if ((13'sd2833/*2833:xpc10*/==xpc10))  xpc10 <= 13'sd2834/*2834:xpc10*/;
                  if ((13'sd2834/*2834:xpc10*/==xpc10))  xpc10 <= 13'sd2835/*2835:xpc10*/;
                  if ((13'sd2835/*2835:xpc10*/==xpc10))  xpc10 <= 13'sd2836/*2836:xpc10*/;
                  if ((13'sd2837/*2837:xpc10*/==xpc10))  xpc10 <= 13'sd2838/*2838:xpc10*/;
                  if ((13'sd2838/*2838:xpc10*/==xpc10))  xpc10 <= 13'sd2839/*2839:xpc10*/;
                  if ((13'sd2839/*2839:xpc10*/==xpc10))  xpc10 <= 13'sd2840/*2840:xpc10*/;
                  if ((13'sd2841/*2841:xpc10*/==xpc10))  xpc10 <= 13'sd2842/*2842:xpc10*/;
                  if ((13'sd2842/*2842:xpc10*/==xpc10))  xpc10 <= 13'sd2843/*2843:xpc10*/;
                  if ((13'sd2843/*2843:xpc10*/==xpc10))  xpc10 <= 13'sd2844/*2844:xpc10*/;
                  if ((13'sd2845/*2845:xpc10*/==xpc10))  xpc10 <= 13'sd2846/*2846:xpc10*/;
                  if ((13'sd2846/*2846:xpc10*/==xpc10))  xpc10 <= 13'sd2847/*2847:xpc10*/;
                  if ((13'sd2847/*2847:xpc10*/==xpc10))  xpc10 <= 13'sd2848/*2848:xpc10*/;
                  if ((13'sd2849/*2849:xpc10*/==xpc10))  xpc10 <= 13'sd2850/*2850:xpc10*/;
                  if ((13'sd2850/*2850:xpc10*/==xpc10))  xpc10 <= 13'sd2851/*2851:xpc10*/;
                  if ((13'sd2851/*2851:xpc10*/==xpc10))  xpc10 <= 13'sd2852/*2852:xpc10*/;
                  if ((13'sd2853/*2853:xpc10*/==xpc10))  xpc10 <= 13'sd2854/*2854:xpc10*/;
                  if ((13'sd2854/*2854:xpc10*/==xpc10))  xpc10 <= 13'sd2855/*2855:xpc10*/;
                  if ((13'sd2855/*2855:xpc10*/==xpc10))  xpc10 <= 13'sd2856/*2856:xpc10*/;
                  if ((13'sd2857/*2857:xpc10*/==xpc10))  xpc10 <= 13'sd2781/*2781:xpc10*/;
                  if ((13'sd2858/*2858:xpc10*/==xpc10))  xpc10 <= 13'sd2859/*2859:xpc10*/;
                  if ((13'sd2859/*2859:xpc10*/==xpc10))  xpc10 <= 13'sd2860/*2860:xpc10*/;
                  if ((13'sd2861/*2861:xpc10*/==xpc10))  xpc10 <= 13'sd2854/*2854:xpc10*/;
                  if ((13'sd2862/*2862:xpc10*/==xpc10))  xpc10 <= 13'sd2863/*2863:xpc10*/;
                  if ((13'sd2863/*2863:xpc10*/==xpc10))  xpc10 <= 13'sd2864/*2864:xpc10*/;
                  if ((13'sd2865/*2865:xpc10*/==xpc10))  xpc10 <= 13'sd2866/*2866:xpc10*/;
                  if ((13'sd2866/*2866:xpc10*/==xpc10))  xpc10 <= 13'sd2867/*2867:xpc10*/;
                  if ((13'sd2867/*2867:xpc10*/==xpc10))  xpc10 <= 13'sd2868/*2868:xpc10*/;
                  if ((13'sd2872/*2872:xpc10*/==xpc10))  xpc10 <= 13'sd2873/*2873:xpc10*/;
                  if ((13'sd2873/*2873:xpc10*/==xpc10))  xpc10 <= 13'sd2874/*2874:xpc10*/;
                  if ((13'sd2874/*2874:xpc10*/==xpc10))  xpc10 <= 13'sd2875/*2875:xpc10*/;
                  if ((13'sd2877/*2877:xpc10*/==xpc10))  xpc10 <= 13'sd2878/*2878:xpc10*/;
                  if ((13'sd2878/*2878:xpc10*/==xpc10))  xpc10 <= 13'sd2879/*2879:xpc10*/;
                  if ((13'sd2879/*2879:xpc10*/==xpc10))  xpc10 <= 13'sd2880/*2880:xpc10*/;
                  if ((13'sd2881/*2881:xpc10*/==xpc10))  xpc10 <= 13'sd2807/*2807:xpc10*/;
                  if ((13'sd2882/*2882:xpc10*/==xpc10))  xpc10 <= 13'sd2883/*2883:xpc10*/;
                  if ((13'sd2883/*2883:xpc10*/==xpc10))  xpc10 <= 13'sd2884/*2884:xpc10*/;
                  if ((13'sd2886/*2886:xpc10*/==xpc10))  xpc10 <= 13'sd2878/*2878:xpc10*/;
                  if ((13'sd2887/*2887:xpc10*/==xpc10))  xpc10 <= 13'sd2888/*2888:xpc10*/;
                  if ((13'sd2888/*2888:xpc10*/==xpc10))  xpc10 <= 13'sd2889/*2889:xpc10*/;
                  if ((13'sd2890/*2890:xpc10*/==xpc10))  xpc10 <= 13'sd2891/*2891:xpc10*/;
                  if ((13'sd2891/*2891:xpc10*/==xpc10))  xpc10 <= 13'sd2892/*2892:xpc10*/;
                  if ((13'sd2892/*2892:xpc10*/==xpc10))  xpc10 <= 13'sd2893/*2893:xpc10*/;
                  if ((13'sd2894/*2894:xpc10*/==xpc10))  xpc10 <= 13'sd2895/*2895:xpc10*/;
                  if ((13'sd2895/*2895:xpc10*/==xpc10))  xpc10 <= 13'sd2896/*2896:xpc10*/;
                  if ((13'sd2896/*2896:xpc10*/==xpc10))  xpc10 <= 13'sd2897/*2897:xpc10*/;
                  if ((13'sd2898/*2898:xpc10*/==xpc10))  xpc10 <= 13'sd2807/*2807:xpc10*/;
                  if ((13'sd2899/*2899:xpc10*/==xpc10))  xpc10 <= 13'sd2900/*2900:xpc10*/;
                  if ((13'sd2900/*2900:xpc10*/==xpc10))  xpc10 <= 13'sd2901/*2901:xpc10*/;
                  if ((13'sd2902/*2902:xpc10*/==xpc10))  xpc10 <= 13'sd2895/*2895:xpc10*/;
                  if ((13'sd2903/*2903:xpc10*/==xpc10))  xpc10 <= 13'sd2904/*2904:xpc10*/;
                  if ((13'sd2904/*2904:xpc10*/==xpc10))  xpc10 <= 13'sd2905/*2905:xpc10*/;
                  if ((13'sd2907/*2907:xpc10*/==xpc10))  xpc10 <= 13'sd2727/*2727:xpc10*/;
                  if ((13'sd2908/*2908:xpc10*/==xpc10))  xpc10 <= 13'sd2909/*2909:xpc10*/;
                  if ((13'sd2909/*2909:xpc10*/==xpc10))  xpc10 <= 13'sd2910/*2910:xpc10*/;
                  if ((13'sd2917/*2917:xpc10*/==xpc10))  xpc10 <= 13'sd2918/*2918:xpc10*/;
                  if ((13'sd2918/*2918:xpc10*/==xpc10))  xpc10 <= 13'sd2919/*2919:xpc10*/;
                  if ((13'sd2919/*2919:xpc10*/==xpc10))  xpc10 <= 13'sd2920/*2920:xpc10*/;
                  if ((13'sd2922/*2922:xpc10*/==xpc10))  xpc10 <= 13'sd2923/*2923:xpc10*/;
                  if ((13'sd2923/*2923:xpc10*/==xpc10))  xpc10 <= 13'sd2924/*2924:xpc10*/;
                  if ((13'sd2924/*2924:xpc10*/==xpc10))  xpc10 <= 13'sd2925/*2925:xpc10*/;
                  if ((13'sd2926/*2926:xpc10*/==xpc10))  xpc10 <= 13'sd2711/*2711:xpc10*/;
                  if ((13'sd2927/*2927:xpc10*/==xpc10))  xpc10 <= 13'sd2928/*2928:xpc10*/;
                  if ((13'sd2928/*2928:xpc10*/==xpc10))  xpc10 <= 13'sd2929/*2929:xpc10*/;
                  if ((13'sd2931/*2931:xpc10*/==xpc10))  xpc10 <= 13'sd2923/*2923:xpc10*/;
                  if ((13'sd2932/*2932:xpc10*/==xpc10))  xpc10 <= 13'sd2933/*2933:xpc10*/;
                  if ((13'sd2933/*2933:xpc10*/==xpc10))  xpc10 <= 13'sd2934/*2934:xpc10*/;
                  if ((13'sd2936/*2936:xpc10*/==xpc10))  xpc10 <= 13'sd2707/*2707:xpc10*/;
                  if ((13'sd2937/*2937:xpc10*/==xpc10))  xpc10 <= 13'sd2938/*2938:xpc10*/;
                  if ((13'sd2938/*2938:xpc10*/==xpc10))  xpc10 <= 13'sd2939/*2939:xpc10*/;
                  if ((13'sd2941/*2941:xpc10*/==xpc10))  xpc10 <= 13'sd2691/*2691:xpc10*/;
                  if ((13'sd2942/*2942:xpc10*/==xpc10))  xpc10 <= 13'sd2943/*2943:xpc10*/;
                  if ((13'sd2943/*2943:xpc10*/==xpc10))  xpc10 <= 13'sd2944/*2944:xpc10*/;
                  if ((13'sd2946/*2946:xpc10*/==xpc10))  xpc10 <= 13'sd2676/*2676:xpc10*/;
                  if ((13'sd2947/*2947:xpc10*/==xpc10))  xpc10 <= 13'sd2948/*2948:xpc10*/;
                  if ((13'sd2948/*2948:xpc10*/==xpc10))  xpc10 <= 13'sd2949/*2949:xpc10*/;
                  if ((13'sd2949/*2949:xpc10*/==xpc10))  xpc10 <= 13'sd2950/*2950:xpc10*/;
                  if ((13'sd2950/*2950:xpc10*/==xpc10))  xpc10 <= 13'sd2663/*2663:xpc10*/;
                  if ((13'sd2951/*2951:xpc10*/==xpc10))  xpc10 <= 13'sd2952/*2952:xpc10*/;
                  if ((13'sd2952/*2952:xpc10*/==xpc10))  xpc10 <= 13'sd2953/*2953:xpc10*/;
                  if ((13'sd2955/*2955:xpc10*/==xpc10))  xpc10 <= 13'sd2956/*2956:xpc10*/;
                  if ((13'sd2956/*2956:xpc10*/==xpc10))  xpc10 <= 13'sd2957/*2957:xpc10*/;
                  if ((13'sd2957/*2957:xpc10*/==xpc10))  xpc10 <= 13'sd2958/*2958:xpc10*/;
                  if ((13'sd2959/*2959:xpc10*/==xpc10))  xpc10 <= 13'sd2960/*2960:xpc10*/;
                  if ((13'sd2960/*2960:xpc10*/==xpc10))  xpc10 <= 13'sd2961/*2961:xpc10*/;
                  if ((13'sd2961/*2961:xpc10*/==xpc10))  xpc10 <= 13'sd2962/*2962:xpc10*/;
                  if ((13'sd2973/*2973:xpc10*/==xpc10))  xpc10 <= 13'sd2974/*2974:xpc10*/;
                  if ((13'sd2974/*2974:xpc10*/==xpc10))  xpc10 <= 13'sd2975/*2975:xpc10*/;
                  if ((13'sd2975/*2975:xpc10*/==xpc10))  xpc10 <= 13'sd2976/*2976:xpc10*/;
                  if ((13'sd2976/*2976:xpc10*/==xpc10))  xpc10 <= 13'sd2977/*2977:xpc10*/;
                  if ((13'sd2977/*2977:xpc10*/==xpc10))  xpc10 <= 13'sd2978/*2978:xpc10*/;
                  if ((13'sd2978/*2978:xpc10*/==xpc10))  xpc10 <= 13'sd2979/*2979:xpc10*/;
                  if ((13'sd2979/*2979:xpc10*/==xpc10))  xpc10 <= 13'sd2980/*2980:xpc10*/;
                  if ((13'sd2980/*2980:xpc10*/==xpc10))  xpc10 <= 13'sd2981/*2981:xpc10*/;
                  if ((13'sd2985/*2985:xpc10*/==xpc10))  xpc10 <= 13'sd2986/*2986:xpc10*/;
                  if ((13'sd2986/*2986:xpc10*/==xpc10))  xpc10 <= 13'sd2987/*2987:xpc10*/;
                  if ((13'sd2987/*2987:xpc10*/==xpc10))  xpc10 <= 13'sd2988/*2988:xpc10*/;
                  if ((13'sd2990/*2990:xpc10*/==xpc10))  xpc10 <= 13'sd2991/*2991:xpc10*/;
                  if ((13'sd2991/*2991:xpc10*/==xpc10))  xpc10 <= 13'sd2992/*2992:xpc10*/;
                  if ((13'sd2992/*2992:xpc10*/==xpc10))  xpc10 <= 13'sd2993/*2993:xpc10*/;
                  if ((13'sd3000/*3000:xpc10*/==xpc10))  xpc10 <= 13'sd3001/*3001:xpc10*/;
                  if ((13'sd3001/*3001:xpc10*/==xpc10))  xpc10 <= 13'sd3002/*3002:xpc10*/;
                  if ((13'sd3002/*3002:xpc10*/==xpc10))  xpc10 <= 13'sd3003/*3003:xpc10*/;
                  if ((13'sd3005/*3005:xpc10*/==xpc10))  xpc10 <= 13'sd3006/*3006:xpc10*/;
                  if ((13'sd3006/*3006:xpc10*/==xpc10))  xpc10 <= 13'sd3007/*3007:xpc10*/;
                  if ((13'sd3007/*3007:xpc10*/==xpc10))  xpc10 <= 13'sd3008/*3008:xpc10*/;
                  if ((13'sd3016/*3016:xpc10*/==xpc10))  xpc10 <= 13'sd3017/*3017:xpc10*/;
                  if ((13'sd3017/*3017:xpc10*/==xpc10))  xpc10 <= 13'sd3018/*3018:xpc10*/;
                  if ((13'sd3018/*3018:xpc10*/==xpc10))  xpc10 <= 13'sd3019/*3019:xpc10*/;
                  if ((13'sd3021/*3021:xpc10*/==xpc10))  xpc10 <= 13'sd3022/*3022:xpc10*/;
                  if ((13'sd3022/*3022:xpc10*/==xpc10))  xpc10 <= 13'sd3023/*3023:xpc10*/;
                  if ((13'sd3023/*3023:xpc10*/==xpc10))  xpc10 <= 13'sd3024/*3024:xpc10*/;
                  if ((13'sd3025/*3025:xpc10*/==xpc10))  xpc10 <= 13'sd3026/*3026:xpc10*/;
                  if ((13'sd3026/*3026:xpc10*/==xpc10))  xpc10 <= 13'sd3027/*3027:xpc10*/;
                  if ((13'sd3027/*3027:xpc10*/==xpc10))  xpc10 <= 13'sd3028/*3028:xpc10*/;
                  if ((13'sd3029/*3029:xpc10*/==xpc10))  xpc10 <= 13'sd3030/*3030:xpc10*/;
                  if ((13'sd3030/*3030:xpc10*/==xpc10))  xpc10 <= 13'sd3031/*3031:xpc10*/;
                  if ((13'sd3031/*3031:xpc10*/==xpc10))  xpc10 <= 13'sd3032/*3032:xpc10*/;
                  if ((13'sd3037/*3037:xpc10*/==xpc10))  xpc10 <= 13'sd3038/*3038:xpc10*/;
                  if ((13'sd3038/*3038:xpc10*/==xpc10))  xpc10 <= 13'sd3039/*3039:xpc10*/;
                  if ((13'sd3039/*3039:xpc10*/==xpc10))  xpc10 <= 13'sd3040/*3040:xpc10*/;
                  if ((13'sd3042/*3042:xpc10*/==xpc10))  xpc10 <= 13'sd3043/*3043:xpc10*/;
                  if ((13'sd3043/*3043:xpc10*/==xpc10))  xpc10 <= 13'sd3044/*3044:xpc10*/;
                  if ((13'sd3044/*3044:xpc10*/==xpc10))  xpc10 <= 13'sd3045/*3045:xpc10*/;
                  if ((13'sd3047/*3047:xpc10*/==xpc10))  xpc10 <= 13'sd2641/*2641:xpc10*/;
                  if ((13'sd3048/*3048:xpc10*/==xpc10))  xpc10 <= 13'sd3049/*3049:xpc10*/;
                  if ((13'sd3049/*3049:xpc10*/==xpc10))  xpc10 <= 13'sd3050/*3050:xpc10*/;
                  if ((13'sd3052/*3052:xpc10*/==xpc10))  xpc10 <= 13'sd3043/*3043:xpc10*/;
                  if ((13'sd3053/*3053:xpc10*/==xpc10))  xpc10 <= 13'sd3054/*3054:xpc10*/;
                  if ((13'sd3054/*3054:xpc10*/==xpc10))  xpc10 <= 13'sd3055/*3055:xpc10*/;
                  if ((13'sd3063/*3063:xpc10*/==xpc10))  xpc10 <= 13'sd3064/*3064:xpc10*/;
                  if ((13'sd3064/*3064:xpc10*/==xpc10))  xpc10 <= 13'sd3065/*3065:xpc10*/;
                  if ((13'sd3065/*3065:xpc10*/==xpc10))  xpc10 <= 13'sd3066/*3066:xpc10*/;
                  if ((13'sd3068/*3068:xpc10*/==xpc10))  xpc10 <= 13'sd3069/*3069:xpc10*/;
                  if ((13'sd3069/*3069:xpc10*/==xpc10))  xpc10 <= 13'sd3070/*3070:xpc10*/;
                  if ((13'sd3070/*3070:xpc10*/==xpc10))  xpc10 <= 13'sd3071/*3071:xpc10*/;
                  if ((13'sd3072/*3072:xpc10*/==xpc10))  xpc10 <= 13'sd3026/*3026:xpc10*/;
                  if ((13'sd3073/*3073:xpc10*/==xpc10))  xpc10 <= 13'sd3074/*3074:xpc10*/;
                  if ((13'sd3074/*3074:xpc10*/==xpc10))  xpc10 <= 13'sd3075/*3075:xpc10*/;
                  if ((13'sd3077/*3077:xpc10*/==xpc10))  xpc10 <= 13'sd3069/*3069:xpc10*/;
                  if ((13'sd3078/*3078:xpc10*/==xpc10))  xpc10 <= 13'sd3079/*3079:xpc10*/;
                  if ((13'sd3079/*3079:xpc10*/==xpc10))  xpc10 <= 13'sd3080/*3080:xpc10*/;
                  if ((13'sd3082/*3082:xpc10*/==xpc10))  xpc10 <= 13'sd3022/*3022:xpc10*/;
                  if ((13'sd3083/*3083:xpc10*/==xpc10))  xpc10 <= 13'sd3084/*3084:xpc10*/;
                  if ((13'sd3084/*3084:xpc10*/==xpc10))  xpc10 <= 13'sd3085/*3085:xpc10*/;
                  if ((13'sd3087/*3087:xpc10*/==xpc10))  xpc10 <= 13'sd3006/*3006:xpc10*/;
                  if ((13'sd3088/*3088:xpc10*/==xpc10))  xpc10 <= 13'sd3089/*3089:xpc10*/;
                  if ((13'sd3089/*3089:xpc10*/==xpc10))  xpc10 <= 13'sd3090/*3090:xpc10*/;
                  if ((13'sd3092/*3092:xpc10*/==xpc10))  xpc10 <= 13'sd2991/*2991:xpc10*/;
                  if ((13'sd3093/*3093:xpc10*/==xpc10))  xpc10 <= 13'sd3094/*3094:xpc10*/;
                  if ((13'sd3094/*3094:xpc10*/==xpc10))  xpc10 <= 13'sd3095/*3095:xpc10*/;
                  if ((13'sd3095/*3095:xpc10*/==xpc10))  xpc10 <= 13'sd3096/*3096:xpc10*/;
                  if ((13'sd3096/*3096:xpc10*/==xpc10))  xpc10 <= 13'sd2978/*2978:xpc10*/;
                  if ((13'sd3097/*3097:xpc10*/==xpc10))  xpc10 <= 13'sd3098/*3098:xpc10*/;
                  if ((13'sd3098/*3098:xpc10*/==xpc10))  xpc10 <= 13'sd3099/*3099:xpc10*/;
                  if ((13'sd3100/*3100:xpc10*/==xpc10))  xpc10 <= 13'sd2960/*2960:xpc10*/;
                  if ((13'sd3101/*3101:xpc10*/==xpc10))  xpc10 <= 13'sd3102/*3102:xpc10*/;
                  if ((13'sd3102/*3102:xpc10*/==xpc10))  xpc10 <= 13'sd3103/*3103:xpc10*/;
                  if ((13'sd3104/*3104:xpc10*/==xpc10))  xpc10 <= 13'sd2593/*2593:xpc10*/;
                  if ((13'sd3105/*3105:xpc10*/==xpc10))  xpc10 <= 13'sd3106/*3106:xpc10*/;
                  if ((13'sd3106/*3106:xpc10*/==xpc10))  xpc10 <= 13'sd3107/*3107:xpc10*/;
                  if ((13'sd3108/*3108:xpc10*/==xpc10))  xpc10 <= 13'sd2531/*2531:xpc10*/;
                  if ((13'sd3109/*3109:xpc10*/==xpc10))  xpc10 <= 13'sd3110/*3110:xpc10*/;
                  if ((13'sd3110/*3110:xpc10*/==xpc10))  xpc10 <= 13'sd3111/*3111:xpc10*/;
                  if ((13'sd3112/*3112:xpc10*/==xpc10))  xpc10 <= 13'sd727/*727:xpc10*/;
                  if ((13'sd3113/*3113:xpc10*/==xpc10))  xpc10 <= 13'sd3114/*3114:xpc10*/;
                  if ((13'sd3114/*3114:xpc10*/==xpc10))  xpc10 <= 13'sd3115/*3115:xpc10*/;
                  if ((13'sd3116/*3116:xpc10*/==xpc10))  xpc10 <= 13'sd716/*716:xpc10*/;
                  if ((13'sd3117/*3117:xpc10*/==xpc10))  xpc10 <= 13'sd3118/*3118:xpc10*/;
                  if ((13'sd3118/*3118:xpc10*/==xpc10))  xpc10 <= 13'sd3119/*3119:xpc10*/;
                  if ((13'sd3121/*3121:xpc10*/==xpc10))  xpc10 <= 13'sd3122/*3122:xpc10*/;
                  if ((13'sd3122/*3122:xpc10*/==xpc10))  xpc10 <= 13'sd3123/*3123:xpc10*/;
                  if ((13'sd3123/*3123:xpc10*/==xpc10))  xpc10 <= 13'sd3124/*3124:xpc10*/;
                  if ((13'sd3125/*3125:xpc10*/==xpc10))  xpc10 <= 13'sd3126/*3126:xpc10*/;
                  if ((13'sd3126/*3126:xpc10*/==xpc10))  xpc10 <= 13'sd3127/*3127:xpc10*/;
                  if ((13'sd3127/*3127:xpc10*/==xpc10))  xpc10 <= 13'sd3128/*3128:xpc10*/;
                  if ((13'sd3132/*3132:xpc10*/==xpc10))  xpc10 <= 13'sd3133/*3133:xpc10*/;
                  if ((13'sd3133/*3133:xpc10*/==xpc10))  xpc10 <= 13'sd3134/*3134:xpc10*/;
                  if ((13'sd3134/*3134:xpc10*/==xpc10))  xpc10 <= 13'sd3135/*3135:xpc10*/;
                  if ((13'sd3137/*3137:xpc10*/==xpc10))  xpc10 <= 13'sd3138/*3138:xpc10*/;
                  if ((13'sd3138/*3138:xpc10*/==xpc10))  xpc10 <= 13'sd3139/*3139:xpc10*/;
                  if ((13'sd3139/*3139:xpc10*/==xpc10))  xpc10 <= 13'sd3140/*3140:xpc10*/;
                  if ((13'sd3141/*3141:xpc10*/==xpc10))  xpc10 <= 13'sd3142/*3142:xpc10*/;
                  if ((13'sd3142/*3142:xpc10*/==xpc10))  xpc10 <= 13'sd3143/*3143:xpc10*/;
                  if ((13'sd3143/*3143:xpc10*/==xpc10))  xpc10 <= 13'sd3144/*3144:xpc10*/;
                  if ((13'sd3146/*3146:xpc10*/==xpc10))  xpc10 <= 13'sd3147/*3147:xpc10*/;
                  if ((13'sd3147/*3147:xpc10*/==xpc10))  xpc10 <= 13'sd3148/*3148:xpc10*/;
                  if ((13'sd3148/*3148:xpc10*/==xpc10))  xpc10 <= 13'sd3149/*3149:xpc10*/;
                  if ((13'sd3153/*3153:xpc10*/==xpc10))  xpc10 <= 13'sd3154/*3154:xpc10*/;
                  if ((13'sd3154/*3154:xpc10*/==xpc10))  xpc10 <= 13'sd3155/*3155:xpc10*/;
                  if ((13'sd3155/*3155:xpc10*/==xpc10))  xpc10 <= 13'sd3156/*3156:xpc10*/;
                  if ((13'sd3157/*3157:xpc10*/==xpc10))  xpc10 <= 13'sd3158/*3158:xpc10*/;
                  if ((13'sd3158/*3158:xpc10*/==xpc10))  xpc10 <= 13'sd3159/*3159:xpc10*/;
                  if ((13'sd3159/*3159:xpc10*/==xpc10))  xpc10 <= 13'sd3160/*3160:xpc10*/;
                  if ((13'sd3161/*3161:xpc10*/==xpc10))  xpc10 <= 13'sd706/*706:xpc10*/;
                  if ((13'sd3162/*3162:xpc10*/==xpc10))  xpc10 <= 13'sd3163/*3163:xpc10*/;
                  if ((13'sd3163/*3163:xpc10*/==xpc10))  xpc10 <= 13'sd3164/*3164:xpc10*/;
                  if ((13'sd3165/*3165:xpc10*/==xpc10))  xpc10 <= 13'sd3158/*3158:xpc10*/;
                  if ((13'sd3166/*3166:xpc10*/==xpc10))  xpc10 <= 13'sd3167/*3167:xpc10*/;
                  if ((13'sd3167/*3167:xpc10*/==xpc10))  xpc10 <= 13'sd3168/*3168:xpc10*/;
                  if ((13'sd3169/*3169:xpc10*/==xpc10))  xpc10 <= 13'sd3126/*3126:xpc10*/;
                  if ((13'sd3170/*3170:xpc10*/==xpc10))  xpc10 <= 13'sd3171/*3171:xpc10*/;
                  if ((13'sd3171/*3171:xpc10*/==xpc10))  xpc10 <= 13'sd3172/*3172:xpc10*/;
                  if ((13'sd3173/*3173:xpc10*/==xpc10))  xpc10 <= 13'sd3174/*3174:xpc10*/;
                  if ((13'sd3174/*3174:xpc10*/==xpc10))  xpc10 <= 13'sd3175/*3175:xpc10*/;
                  if ((13'sd3175/*3175:xpc10*/==xpc10))  xpc10 <= 13'sd3176/*3176:xpc10*/;
                  if ((13'sd3177/*3177:xpc10*/==xpc10))  xpc10 <= 13'sd694/*694:xpc10*/;
                  if ((13'sd3178/*3178:xpc10*/==xpc10))  xpc10 <= 13'sd3179/*3179:xpc10*/;
                  if ((13'sd3179/*3179:xpc10*/==xpc10))  xpc10 <= 13'sd3180/*3180:xpc10*/;
                  if ((13'sd3181/*3181:xpc10*/==xpc10))  xpc10 <= 13'sd3182/*3182:xpc10*/;
                  if ((13'sd3182/*3182:xpc10*/==xpc10))  xpc10 <= 13'sd3183/*3183:xpc10*/;
                  if ((13'sd3183/*3183:xpc10*/==xpc10))  xpc10 <= 13'sd3184/*3184:xpc10*/;
                  if ((13'sd3185/*3185:xpc10*/==xpc10))  xpc10 <= 13'sd694/*694:xpc10*/;
                  if ((13'sd3186/*3186:xpc10*/==xpc10))  xpc10 <= 13'sd3187/*3187:xpc10*/;
                  if ((13'sd3187/*3187:xpc10*/==xpc10))  xpc10 <= 13'sd3188/*3188:xpc10*/;
                  if ((13'sd3189/*3189:xpc10*/==xpc10))  xpc10 <= 13'sd694/*694:xpc10*/;
                  if ((13'sd3190/*3190:xpc10*/==xpc10))  xpc10 <= 13'sd3191/*3191:xpc10*/;
                  if ((13'sd3191/*3191:xpc10*/==xpc10))  xpc10 <= 13'sd3192/*3192:xpc10*/;
                  if ((13'sd3193/*3193:xpc10*/==xpc10))  xpc10 <= 13'sd675/*675:xpc10*/;
                  if ((13'sd3194/*3194:xpc10*/==xpc10))  xpc10 <= 13'sd3195/*3195:xpc10*/;
                  if ((13'sd3195/*3195:xpc10*/==xpc10))  xpc10 <= 13'sd3196/*3196:xpc10*/;
                  if ((13'sd3197/*3197:xpc10*/==xpc10))  xpc10 <= 13'sd665/*665:xpc10*/;
                  if ((13'sd3198/*3198:xpc10*/==xpc10))  xpc10 <= 13'sd3199/*3199:xpc10*/;
                  if ((13'sd3199/*3199:xpc10*/==xpc10))  xpc10 <= 13'sd3200/*3200:xpc10*/;
                  if ((13'sd3201/*3201:xpc10*/==xpc10))  xpc10 <= 13'sd3202/*3202:xpc10*/;
                  if ((13'sd3202/*3202:xpc10*/==xpc10))  xpc10 <= 13'sd3203/*3203:xpc10*/;
                  if ((13'sd3203/*3203:xpc10*/==xpc10))  xpc10 <= 13'sd3204/*3204:xpc10*/;
                  if ((13'sd3205/*3205:xpc10*/==xpc10))  xpc10 <= 13'sd3206/*3206:xpc10*/;
                  if ((13'sd3206/*3206:xpc10*/==xpc10))  xpc10 <= 13'sd3207/*3207:xpc10*/;
                  if ((13'sd3207/*3207:xpc10*/==xpc10))  xpc10 <= 13'sd3208/*3208:xpc10*/;
                  if ((13'sd3208/*3208:xpc10*/==xpc10))  xpc10 <= 13'sd3209/*3209:xpc10*/;
                  if ((13'sd3210/*3210:xpc10*/==xpc10))  xpc10 <= 13'sd698/*698:xpc10*/;
                  if ((13'sd3211/*3211:xpc10*/==xpc10))  xpc10 <= 13'sd3212/*3212:xpc10*/;
                  if ((13'sd3212/*3212:xpc10*/==xpc10))  xpc10 <= 13'sd3213/*3213:xpc10*/;
                  if ((13'sd3214/*3214:xpc10*/==xpc10))  xpc10 <= 13'sd3215/*3215:xpc10*/;
                  if ((13'sd3215/*3215:xpc10*/==xpc10))  xpc10 <= 13'sd3216/*3216:xpc10*/;
                  if ((13'sd3216/*3216:xpc10*/==xpc10))  xpc10 <= 13'sd3217/*3217:xpc10*/;
                  if ((13'sd3218/*3218:xpc10*/==xpc10))  xpc10 <= 13'sd3219/*3219:xpc10*/;
                  if ((13'sd3219/*3219:xpc10*/==xpc10))  xpc10 <= 13'sd3220/*3220:xpc10*/;
                  if ((13'sd3220/*3220:xpc10*/==xpc10))  xpc10 <= 13'sd3221/*3221:xpc10*/;
                  if ((13'sd3222/*3222:xpc10*/==xpc10))  xpc10 <= 13'sd698/*698:xpc10*/;
                  if ((13'sd3223/*3223:xpc10*/==xpc10))  xpc10 <= 13'sd3224/*3224:xpc10*/;
                  if ((13'sd3224/*3224:xpc10*/==xpc10))  xpc10 <= 13'sd3225/*3225:xpc10*/;
                  if ((13'sd3226/*3226:xpc10*/==xpc10))  xpc10 <= 13'sd3219/*3219:xpc10*/;
                  if ((13'sd3227/*3227:xpc10*/==xpc10))  xpc10 <= 13'sd3228/*3228:xpc10*/;
                  if ((13'sd3228/*3228:xpc10*/==xpc10))  xpc10 <= 13'sd3229/*3229:xpc10*/;
                  if ((13'sd3230/*3230:xpc10*/==xpc10))  xpc10 <= 13'sd3231/*3231:xpc10*/;
                  if ((13'sd3231/*3231:xpc10*/==xpc10))  xpc10 <= 13'sd3232/*3232:xpc10*/;
                  if ((13'sd3232/*3232:xpc10*/==xpc10))  xpc10 <= 13'sd3233/*3233:xpc10*/;
                  if ((13'sd3234/*3234:xpc10*/==xpc10))  xpc10 <= 13'sd3235/*3235:xpc10*/;
                  if ((13'sd3235/*3235:xpc10*/==xpc10))  xpc10 <= 13'sd3236/*3236:xpc10*/;
                  if ((13'sd3236/*3236:xpc10*/==xpc10))  xpc10 <= 13'sd3237/*3237:xpc10*/;
                  if ((13'sd3240/*3240:xpc10*/==xpc10))  xpc10 <= 13'sd3241/*3241:xpc10*/;
                  if ((13'sd3241/*3241:xpc10*/==xpc10))  xpc10 <= 13'sd3242/*3242:xpc10*/;
                  if ((13'sd3242/*3242:xpc10*/==xpc10))  xpc10 <= 13'sd3243/*3243:xpc10*/;
                  if ((13'sd3244/*3244:xpc10*/==xpc10))  xpc10 <= 13'sd3245/*3245:xpc10*/;
                  if ((13'sd3245/*3245:xpc10*/==xpc10))  xpc10 <= 13'sd3246/*3246:xpc10*/;
                  if ((13'sd3246/*3246:xpc10*/==xpc10))  xpc10 <= 13'sd3247/*3247:xpc10*/;
                  if ((13'sd3250/*3250:xpc10*/==xpc10))  xpc10 <= 13'sd3251/*3251:xpc10*/;
                  if ((13'sd3251/*3251:xpc10*/==xpc10))  xpc10 <= 13'sd3252/*3252:xpc10*/;
                  if ((13'sd3252/*3252:xpc10*/==xpc10))  xpc10 <= 13'sd3253/*3253:xpc10*/;
                  if ((13'sd3254/*3254:xpc10*/==xpc10))  xpc10 <= 13'sd3255/*3255:xpc10*/;
                  if ((13'sd3255/*3255:xpc10*/==xpc10))  xpc10 <= 13'sd3256/*3256:xpc10*/;
                  if ((13'sd3256/*3256:xpc10*/==xpc10))  xpc10 <= 13'sd3257/*3257:xpc10*/;
                  if ((13'sd3261/*3261:xpc10*/==xpc10))  xpc10 <= 13'sd3262/*3262:xpc10*/;
                  if ((13'sd3262/*3262:xpc10*/==xpc10))  xpc10 <= 13'sd3263/*3263:xpc10*/;
                  if ((13'sd3263/*3263:xpc10*/==xpc10))  xpc10 <= 13'sd3264/*3264:xpc10*/;
                  if ((13'sd3264/*3264:xpc10*/==xpc10))  xpc10 <= 13'sd3265/*3265:xpc10*/;
                  if ((13'sd3265/*3265:xpc10*/==xpc10))  xpc10 <= 13'sd3266/*3266:xpc10*/;
                  if ((13'sd3266/*3266:xpc10*/==xpc10))  xpc10 <= 13'sd3267/*3267:xpc10*/;
                  if ((13'sd3267/*3267:xpc10*/==xpc10))  xpc10 <= 13'sd3268/*3268:xpc10*/;
                  if ((13'sd3269/*3269:xpc10*/==xpc10))  xpc10 <= 13'sd3270/*3270:xpc10*/;
                  if ((13'sd3270/*3270:xpc10*/==xpc10))  xpc10 <= 13'sd3271/*3271:xpc10*/;
                  if ((13'sd3271/*3271:xpc10*/==xpc10))  xpc10 <= 13'sd3272/*3272:xpc10*/;
                  if ((13'sd3273/*3273:xpc10*/==xpc10))  xpc10 <= 13'sd3274/*3274:xpc10*/;
                  if ((13'sd3274/*3274:xpc10*/==xpc10))  xpc10 <= 13'sd3275/*3275:xpc10*/;
                  if ((13'sd3275/*3275:xpc10*/==xpc10))  xpc10 <= 13'sd3276/*3276:xpc10*/;
                  if ((13'sd3277/*3277:xpc10*/==xpc10))  xpc10 <= 13'sd698/*698:xpc10*/;
                  if ((13'sd3278/*3278:xpc10*/==xpc10))  xpc10 <= 13'sd3279/*3279:xpc10*/;
                  if ((13'sd3279/*3279:xpc10*/==xpc10))  xpc10 <= 13'sd3280/*3280:xpc10*/;
                  if ((13'sd3281/*3281:xpc10*/==xpc10))  xpc10 <= 13'sd3282/*3282:xpc10*/;
                  if ((13'sd3282/*3282:xpc10*/==xpc10))  xpc10 <= 13'sd3283/*3283:xpc10*/;
                  if ((13'sd3283/*3283:xpc10*/==xpc10))  xpc10 <= 13'sd3284/*3284:xpc10*/;
                  if ((13'sd3285/*3285:xpc10*/==xpc10))  xpc10 <= 13'sd3274/*3274:xpc10*/;
                  if ((13'sd3286/*3286:xpc10*/==xpc10))  xpc10 <= 13'sd3287/*3287:xpc10*/;
                  if ((13'sd3287/*3287:xpc10*/==xpc10))  xpc10 <= 13'sd3288/*3288:xpc10*/;
                  if ((13'sd3289/*3289:xpc10*/==xpc10))  xpc10 <= 13'sd3290/*3290:xpc10*/;
                  if ((13'sd3290/*3290:xpc10*/==xpc10))  xpc10 <= 13'sd3291/*3291:xpc10*/;
                  if ((13'sd3291/*3291:xpc10*/==xpc10))  xpc10 <= 13'sd3292/*3292:xpc10*/;
                  if ((13'sd3293/*3293:xpc10*/==xpc10))  xpc10 <= 13'sd3274/*3274:xpc10*/;
                  if ((13'sd3294/*3294:xpc10*/==xpc10))  xpc10 <= 13'sd3295/*3295:xpc10*/;
                  if ((13'sd3295/*3295:xpc10*/==xpc10))  xpc10 <= 13'sd3296/*3296:xpc10*/;
                  if ((13'sd3297/*3297:xpc10*/==xpc10))  xpc10 <= 13'sd3274/*3274:xpc10*/;
                  if ((13'sd3298/*3298:xpc10*/==xpc10))  xpc10 <= 13'sd3299/*3299:xpc10*/;
                  if ((13'sd3299/*3299:xpc10*/==xpc10))  xpc10 <= 13'sd3300/*3300:xpc10*/;
                  if ((13'sd3301/*3301:xpc10*/==xpc10))  xpc10 <= 13'sd3255/*3255:xpc10*/;
                  if ((13'sd3302/*3302:xpc10*/==xpc10))  xpc10 <= 13'sd3303/*3303:xpc10*/;
                  if ((13'sd3303/*3303:xpc10*/==xpc10))  xpc10 <= 13'sd3304/*3304:xpc10*/;
                  if ((13'sd3305/*3305:xpc10*/==xpc10))  xpc10 <= 13'sd3245/*3245:xpc10*/;
                  if ((13'sd3306/*3306:xpc10*/==xpc10))  xpc10 <= 13'sd3307/*3307:xpc10*/;
                  if ((13'sd3307/*3307:xpc10*/==xpc10))  xpc10 <= 13'sd3308/*3308:xpc10*/;
                  if ((13'sd3309/*3309:xpc10*/==xpc10))  xpc10 <= 13'sd3310/*3310:xpc10*/;
                  if ((13'sd3310/*3310:xpc10*/==xpc10))  xpc10 <= 13'sd3311/*3311:xpc10*/;
                  if ((13'sd3311/*3311:xpc10*/==xpc10))  xpc10 <= 13'sd3312/*3312:xpc10*/;
                  if ((13'sd3313/*3313:xpc10*/==xpc10))  xpc10 <= 13'sd3314/*3314:xpc10*/;
                  if ((13'sd3314/*3314:xpc10*/==xpc10))  xpc10 <= 13'sd3315/*3315:xpc10*/;
                  if ((13'sd3315/*3315:xpc10*/==xpc10))  xpc10 <= 13'sd3316/*3316:xpc10*/;
                  if ((13'sd3316/*3316:xpc10*/==xpc10))  xpc10 <= 13'sd3317/*3317:xpc10*/;
                  if ((13'sd3318/*3318:xpc10*/==xpc10))  xpc10 <= 13'sd698/*698:xpc10*/;
                  if ((13'sd3319/*3319:xpc10*/==xpc10))  xpc10 <= 13'sd3320/*3320:xpc10*/;
                  if ((13'sd3320/*3320:xpc10*/==xpc10))  xpc10 <= 13'sd3321/*3321:xpc10*/;
                  if ((13'sd3322/*3322:xpc10*/==xpc10))  xpc10 <= 13'sd3323/*3323:xpc10*/;
                  if ((13'sd3323/*3323:xpc10*/==xpc10))  xpc10 <= 13'sd3324/*3324:xpc10*/;
                  if ((13'sd3324/*3324:xpc10*/==xpc10))  xpc10 <= 13'sd3325/*3325:xpc10*/;
                  if ((13'sd3326/*3326:xpc10*/==xpc10))  xpc10 <= 13'sd3327/*3327:xpc10*/;
                  if ((13'sd3327/*3327:xpc10*/==xpc10))  xpc10 <= 13'sd3328/*3328:xpc10*/;
                  if ((13'sd3328/*3328:xpc10*/==xpc10))  xpc10 <= 13'sd3329/*3329:xpc10*/;
                  if ((13'sd3330/*3330:xpc10*/==xpc10))  xpc10 <= 13'sd698/*698:xpc10*/;
                  if ((13'sd3331/*3331:xpc10*/==xpc10))  xpc10 <= 13'sd3332/*3332:xpc10*/;
                  if ((13'sd3332/*3332:xpc10*/==xpc10))  xpc10 <= 13'sd3333/*3333:xpc10*/;
                  if ((13'sd3334/*3334:xpc10*/==xpc10))  xpc10 <= 13'sd3327/*3327:xpc10*/;
                  if ((13'sd3335/*3335:xpc10*/==xpc10))  xpc10 <= 13'sd3336/*3336:xpc10*/;
                  if ((13'sd3336/*3336:xpc10*/==xpc10))  xpc10 <= 13'sd3337/*3337:xpc10*/;
                  if ((13'sd3338/*3338:xpc10*/==xpc10))  xpc10 <= 13'sd3339/*3339:xpc10*/;
                  if ((13'sd3339/*3339:xpc10*/==xpc10))  xpc10 <= 13'sd3340/*3340:xpc10*/;
                  if ((13'sd3340/*3340:xpc10*/==xpc10))  xpc10 <= 13'sd3341/*3341:xpc10*/;
                  if ((13'sd3342/*3342:xpc10*/==xpc10))  xpc10 <= 13'sd3343/*3343:xpc10*/;
                  if ((13'sd3343/*3343:xpc10*/==xpc10))  xpc10 <= 13'sd3344/*3344:xpc10*/;
                  if ((13'sd3344/*3344:xpc10*/==xpc10))  xpc10 <= 13'sd3345/*3345:xpc10*/;
                  if ((13'sd3346/*3346:xpc10*/==xpc10))  xpc10 <= 13'sd3347/*3347:xpc10*/;
                  if ((13'sd3347/*3347:xpc10*/==xpc10))  xpc10 <= 13'sd3348/*3348:xpc10*/;
                  if ((13'sd3348/*3348:xpc10*/==xpc10))  xpc10 <= 13'sd3349/*3349:xpc10*/;
                  if ((13'sd3350/*3350:xpc10*/==xpc10))  xpc10 <= 13'sd3351/*3351:xpc10*/;
                  if ((13'sd3351/*3351:xpc10*/==xpc10))  xpc10 <= 13'sd3352/*3352:xpc10*/;
                  if ((13'sd3352/*3352:xpc10*/==xpc10))  xpc10 <= 13'sd3353/*3353:xpc10*/;
                  if ((13'sd3354/*3354:xpc10*/==xpc10))  xpc10 <= 13'sd698/*698:xpc10*/;
                  if ((13'sd3355/*3355:xpc10*/==xpc10))  xpc10 <= 13'sd3356/*3356:xpc10*/;
                  if ((13'sd3356/*3356:xpc10*/==xpc10))  xpc10 <= 13'sd3357/*3357:xpc10*/;
                  if ((13'sd3358/*3358:xpc10*/==xpc10))  xpc10 <= 13'sd3351/*3351:xpc10*/;
                  if ((13'sd3359/*3359:xpc10*/==xpc10))  xpc10 <= 13'sd3360/*3360:xpc10*/;
                  if ((13'sd3360/*3360:xpc10*/==xpc10))  xpc10 <= 13'sd3361/*3361:xpc10*/;
                  if ((13'sd3364/*3364:xpc10*/==xpc10))  xpc10 <= 13'sd3365/*3365:xpc10*/;
                  if ((13'sd3365/*3365:xpc10*/==xpc10))  xpc10 <= 13'sd3366/*3366:xpc10*/;
                  if ((13'sd3366/*3366:xpc10*/==xpc10))  xpc10 <= 13'sd3367/*3367:xpc10*/;
                  if ((13'sd3368/*3368:xpc10*/==xpc10))  xpc10 <= 13'sd3369/*3369:xpc10*/;
                  if ((13'sd3369/*3369:xpc10*/==xpc10))  xpc10 <= 13'sd3370/*3370:xpc10*/;
                  if ((13'sd3370/*3370:xpc10*/==xpc10))  xpc10 <= 13'sd3371/*3371:xpc10*/;
                  if ((13'sd3374/*3374:xpc10*/==xpc10))  xpc10 <= 13'sd3375/*3375:xpc10*/;
                  if ((13'sd3375/*3375:xpc10*/==xpc10))  xpc10 <= 13'sd3376/*3376:xpc10*/;
                  if ((13'sd3376/*3376:xpc10*/==xpc10))  xpc10 <= 13'sd3377/*3377:xpc10*/;
                  if ((13'sd3379/*3379:xpc10*/==xpc10))  xpc10 <= 13'sd3380/*3380:xpc10*/;
                  if ((13'sd3380/*3380:xpc10*/==xpc10))  xpc10 <= 13'sd3381/*3381:xpc10*/;
                  if ((13'sd3381/*3381:xpc10*/==xpc10))  xpc10 <= 13'sd3382/*3382:xpc10*/;
                  if ((13'sd3383/*3383:xpc10*/==xpc10))  xpc10 <= 13'sd3384/*3384:xpc10*/;
                  if ((13'sd3384/*3384:xpc10*/==xpc10))  xpc10 <= 13'sd3385/*3385:xpc10*/;
                  if ((13'sd3385/*3385:xpc10*/==xpc10))  xpc10 <= 13'sd3386/*3386:xpc10*/;
                  if ((13'sd3388/*3388:xpc10*/==xpc10))  xpc10 <= 13'sd3389/*3389:xpc10*/;
                  if ((13'sd3389/*3389:xpc10*/==xpc10))  xpc10 <= 13'sd3390/*3390:xpc10*/;
                  if ((13'sd3390/*3390:xpc10*/==xpc10))  xpc10 <= 13'sd3391/*3391:xpc10*/;
                  if ((13'sd3396/*3396:xpc10*/==xpc10))  xpc10 <= 13'sd3397/*3397:xpc10*/;
                  if ((13'sd3397/*3397:xpc10*/==xpc10))  xpc10 <= 13'sd3398/*3398:xpc10*/;
                  if ((13'sd3398/*3398:xpc10*/==xpc10))  xpc10 <= 13'sd3399/*3399:xpc10*/;
                  if ((13'sd3400/*3400:xpc10*/==xpc10))  xpc10 <= 13'sd3401/*3401:xpc10*/;
                  if ((13'sd3401/*3401:xpc10*/==xpc10))  xpc10 <= 13'sd3402/*3402:xpc10*/;
                  if ((13'sd3402/*3402:xpc10*/==xpc10))  xpc10 <= 13'sd3403/*3403:xpc10*/;
                  if ((13'sd3404/*3404:xpc10*/==xpc10))  xpc10 <= 13'sd3405/*3405:xpc10*/;
                  if ((13'sd3405/*3405:xpc10*/==xpc10))  xpc10 <= 13'sd3406/*3406:xpc10*/;
                  if ((13'sd3406/*3406:xpc10*/==xpc10))  xpc10 <= 13'sd3407/*3407:xpc10*/;
                  if ((13'sd3408/*3408:xpc10*/==xpc10))  xpc10 <= 13'sd3409/*3409:xpc10*/;
                  if ((13'sd3409/*3409:xpc10*/==xpc10))  xpc10 <= 13'sd3410/*3410:xpc10*/;
                  if ((13'sd3410/*3410:xpc10*/==xpc10))  xpc10 <= 13'sd3411/*3411:xpc10*/;
                  if ((13'sd3412/*3412:xpc10*/==xpc10))  xpc10 <= 13'sd3413/*3413:xpc10*/;
                  if ((13'sd3413/*3413:xpc10*/==xpc10))  xpc10 <= 13'sd3414/*3414:xpc10*/;
                  if ((13'sd3414/*3414:xpc10*/==xpc10))  xpc10 <= 13'sd3415/*3415:xpc10*/;
                  if ((13'sd3416/*3416:xpc10*/==xpc10))  xpc10 <= 13'sd698/*698:xpc10*/;
                  if ((13'sd3417/*3417:xpc10*/==xpc10))  xpc10 <= 13'sd3418/*3418:xpc10*/;
                  if ((13'sd3418/*3418:xpc10*/==xpc10))  xpc10 <= 13'sd3419/*3419:xpc10*/;
                  if ((13'sd3420/*3420:xpc10*/==xpc10))  xpc10 <= 13'sd3413/*3413:xpc10*/;
                  if ((13'sd3421/*3421:xpc10*/==xpc10))  xpc10 <= 13'sd3422/*3422:xpc10*/;
                  if ((13'sd3422/*3422:xpc10*/==xpc10))  xpc10 <= 13'sd3423/*3423:xpc10*/;
                  if ((13'sd3426/*3426:xpc10*/==xpc10))  xpc10 <= 13'sd3427/*3427:xpc10*/;
                  if ((13'sd3427/*3427:xpc10*/==xpc10))  xpc10 <= 13'sd3428/*3428:xpc10*/;
                  if ((13'sd3428/*3428:xpc10*/==xpc10))  xpc10 <= 13'sd3429/*3429:xpc10*/;
                  if ((13'sd3430/*3430:xpc10*/==xpc10))  xpc10 <= 13'sd3431/*3431:xpc10*/;
                  if ((13'sd3431/*3431:xpc10*/==xpc10))  xpc10 <= 13'sd3432/*3432:xpc10*/;
                  if ((13'sd3432/*3432:xpc10*/==xpc10))  xpc10 <= 13'sd3433/*3433:xpc10*/;
                  if ((13'sd3436/*3436:xpc10*/==xpc10))  xpc10 <= 13'sd3437/*3437:xpc10*/;
                  if ((13'sd3437/*3437:xpc10*/==xpc10))  xpc10 <= 13'sd3438/*3438:xpc10*/;
                  if ((13'sd3438/*3438:xpc10*/==xpc10))  xpc10 <= 13'sd3439/*3439:xpc10*/;
                  if ((13'sd3441/*3441:xpc10*/==xpc10))  xpc10 <= 13'sd3442/*3442:xpc10*/;
                  if ((13'sd3442/*3442:xpc10*/==xpc10))  xpc10 <= 13'sd3443/*3443:xpc10*/;
                  if ((13'sd3443/*3443:xpc10*/==xpc10))  xpc10 <= 13'sd3444/*3444:xpc10*/;
                  if ((13'sd3445/*3445:xpc10*/==xpc10))  xpc10 <= 13'sd3446/*3446:xpc10*/;
                  if ((13'sd3446/*3446:xpc10*/==xpc10))  xpc10 <= 13'sd3447/*3447:xpc10*/;
                  if ((13'sd3447/*3447:xpc10*/==xpc10))  xpc10 <= 13'sd3448/*3448:xpc10*/;
                  if ((13'sd3450/*3450:xpc10*/==xpc10))  xpc10 <= 13'sd3451/*3451:xpc10*/;
                  if ((13'sd3451/*3451:xpc10*/==xpc10))  xpc10 <= 13'sd3452/*3452:xpc10*/;
                  if ((13'sd3452/*3452:xpc10*/==xpc10))  xpc10 <= 13'sd3453/*3453:xpc10*/;
                  if ((13'sd3458/*3458:xpc10*/==xpc10))  xpc10 <= 13'sd3459/*3459:xpc10*/;
                  if ((13'sd3459/*3459:xpc10*/==xpc10))  xpc10 <= 13'sd3460/*3460:xpc10*/;
                  if ((13'sd3460/*3460:xpc10*/==xpc10))  xpc10 <= 13'sd3461/*3461:xpc10*/;
                  if ((13'sd3474/*3474:xpc10*/==xpc10))  xpc10 <= 13'sd3475/*3475:xpc10*/;
                  if ((13'sd3475/*3475:xpc10*/==xpc10))  xpc10 <= 13'sd3476/*3476:xpc10*/;
                  if ((13'sd3476/*3476:xpc10*/==xpc10))  xpc10 <= 13'sd3477/*3477:xpc10*/;
                  if ((13'sd3477/*3477:xpc10*/==xpc10))  xpc10 <= 13'sd3478/*3478:xpc10*/;
                  if ((13'sd3478/*3478:xpc10*/==xpc10))  xpc10 <= 13'sd3479/*3479:xpc10*/;
                  if ((13'sd3479/*3479:xpc10*/==xpc10))  xpc10 <= 13'sd3480/*3480:xpc10*/;
                  if ((13'sd3480/*3480:xpc10*/==xpc10))  xpc10 <= 13'sd3481/*3481:xpc10*/;
                  if ((13'sd3481/*3481:xpc10*/==xpc10))  xpc10 <= 13'sd3482/*3482:xpc10*/;
                  if ((13'sd3486/*3486:xpc10*/==xpc10))  xpc10 <= 13'sd3487/*3487:xpc10*/;
                  if ((13'sd3487/*3487:xpc10*/==xpc10))  xpc10 <= 13'sd3488/*3488:xpc10*/;
                  if ((13'sd3488/*3488:xpc10*/==xpc10))  xpc10 <= 13'sd3489/*3489:xpc10*/;
                  if ((13'sd3491/*3491:xpc10*/==xpc10))  xpc10 <= 13'sd3492/*3492:xpc10*/;
                  if ((13'sd3492/*3492:xpc10*/==xpc10))  xpc10 <= 13'sd3493/*3493:xpc10*/;
                  if ((13'sd3493/*3493:xpc10*/==xpc10))  xpc10 <= 13'sd3494/*3494:xpc10*/;
                  if ((13'sd3501/*3501:xpc10*/==xpc10))  xpc10 <= 13'sd3502/*3502:xpc10*/;
                  if ((13'sd3502/*3502:xpc10*/==xpc10))  xpc10 <= 13'sd3503/*3503:xpc10*/;
                  if ((13'sd3503/*3503:xpc10*/==xpc10))  xpc10 <= 13'sd3504/*3504:xpc10*/;
                  if ((13'sd3506/*3506:xpc10*/==xpc10))  xpc10 <= 13'sd3507/*3507:xpc10*/;
                  if ((13'sd3507/*3507:xpc10*/==xpc10))  xpc10 <= 13'sd3508/*3508:xpc10*/;
                  if ((13'sd3508/*3508:xpc10*/==xpc10))  xpc10 <= 13'sd3509/*3509:xpc10*/;
                  if ((13'sd3516/*3516:xpc10*/==xpc10))  xpc10 <= 13'sd3517/*3517:xpc10*/;
                  if ((13'sd3517/*3517:xpc10*/==xpc10))  xpc10 <= 13'sd3518/*3518:xpc10*/;
                  if ((13'sd3518/*3518:xpc10*/==xpc10))  xpc10 <= 13'sd3519/*3519:xpc10*/;
                  if ((13'sd3521/*3521:xpc10*/==xpc10))  xpc10 <= 13'sd3522/*3522:xpc10*/;
                  if ((13'sd3522/*3522:xpc10*/==xpc10))  xpc10 <= 13'sd3523/*3523:xpc10*/;
                  if ((13'sd3523/*3523:xpc10*/==xpc10))  xpc10 <= 13'sd3524/*3524:xpc10*/;
                  if ((13'sd3526/*3526:xpc10*/==xpc10))  xpc10 <= 13'sd3527/*3527:xpc10*/;
                  if ((13'sd3527/*3527:xpc10*/==xpc10))  xpc10 <= 13'sd3528/*3528:xpc10*/;
                  if ((13'sd3528/*3528:xpc10*/==xpc10))  xpc10 <= 13'sd3529/*3529:xpc10*/;
                  if ((13'sd3531/*3531:xpc10*/==xpc10))  xpc10 <= 13'sd3532/*3532:xpc10*/;
                  if ((13'sd3532/*3532:xpc10*/==xpc10))  xpc10 <= 13'sd3533/*3533:xpc10*/;
                  if ((13'sd3533/*3533:xpc10*/==xpc10))  xpc10 <= 13'sd3534/*3534:xpc10*/;
                  if ((13'sd3536/*3536:xpc10*/==xpc10))  xpc10 <= 13'sd3537/*3537:xpc10*/;
                  if ((13'sd3537/*3537:xpc10*/==xpc10))  xpc10 <= 13'sd3538/*3538:xpc10*/;
                  if ((13'sd3539/*3539:xpc10*/==xpc10))  xpc10 <= 13'sd3540/*3540:xpc10*/;
                  if ((13'sd3540/*3540:xpc10*/==xpc10))  xpc10 <= 13'sd3541/*3541:xpc10*/;
                  if ((13'sd3541/*3541:xpc10*/==xpc10))  xpc10 <= 13'sd3542/*3542:xpc10*/;
                  if ((13'sd3544/*3544:xpc10*/==xpc10))  xpc10 <= 13'sd3545/*3545:xpc10*/;
                  if ((13'sd3545/*3545:xpc10*/==xpc10))  xpc10 <= 13'sd3546/*3546:xpc10*/;
                  if ((13'sd3546/*3546:xpc10*/==xpc10))  xpc10 <= 13'sd3547/*3547:xpc10*/;
                  if ((13'sd3548/*3548:xpc10*/==xpc10))  xpc10 <= 13'sd3549/*3549:xpc10*/;
                  if ((13'sd3549/*3549:xpc10*/==xpc10))  xpc10 <= 13'sd3550/*3550:xpc10*/;
                  if ((13'sd3550/*3550:xpc10*/==xpc10))  xpc10 <= 13'sd3551/*3551:xpc10*/;
                  if ((13'sd3552/*3552:xpc10*/==xpc10))  xpc10 <= 13'sd3553/*3553:xpc10*/;
                  if ((13'sd3553/*3553:xpc10*/==xpc10))  xpc10 <= 13'sd3554/*3554:xpc10*/;
                  if ((13'sd3554/*3554:xpc10*/==xpc10))  xpc10 <= 13'sd3555/*3555:xpc10*/;
                  if ((13'sd3556/*3556:xpc10*/==xpc10))  xpc10 <= 13'sd3557/*3557:xpc10*/;
                  if ((13'sd3557/*3557:xpc10*/==xpc10))  xpc10 <= 13'sd3558/*3558:xpc10*/;
                  if ((13'sd3558/*3558:xpc10*/==xpc10))  xpc10 <= 13'sd3559/*3559:xpc10*/;
                  if ((13'sd3559/*3559:xpc10*/==xpc10))  xpc10 <= 13'sd3560/*3560:xpc10*/;
                  if ((13'sd3561/*3561:xpc10*/==xpc10))  xpc10 <= 13'sd3562/*3562:xpc10*/;
                  if ((13'sd3562/*3562:xpc10*/==xpc10))  xpc10 <= 13'sd3563/*3563:xpc10*/;
                  if ((13'sd3563/*3563:xpc10*/==xpc10))  xpc10 <= 13'sd3564/*3564:xpc10*/;
                  if ((13'sd3565/*3565:xpc10*/==xpc10))  xpc10 <= 13'sd3566/*3566:xpc10*/;
                  if ((13'sd3566/*3566:xpc10*/==xpc10))  xpc10 <= 13'sd3567/*3567:xpc10*/;
                  if ((13'sd3567/*3567:xpc10*/==xpc10))  xpc10 <= 13'sd3568/*3568:xpc10*/;
                  if ((13'sd3572/*3572:xpc10*/==xpc10))  xpc10 <= 13'sd3573/*3573:xpc10*/;
                  if ((13'sd3573/*3573:xpc10*/==xpc10))  xpc10 <= 13'sd3574/*3574:xpc10*/;
                  if ((13'sd3574/*3574:xpc10*/==xpc10))  xpc10 <= 13'sd3575/*3575:xpc10*/;
                  if ((13'sd3577/*3577:xpc10*/==xpc10))  xpc10 <= 13'sd3578/*3578:xpc10*/;
                  if ((13'sd3578/*3578:xpc10*/==xpc10))  xpc10 <= 13'sd3579/*3579:xpc10*/;
                  if ((13'sd3579/*3579:xpc10*/==xpc10))  xpc10 <= 13'sd3580/*3580:xpc10*/;
                  if ((13'sd3581/*3581:xpc10*/==xpc10))  xpc10 <= 13'sd3582/*3582:xpc10*/;
                  if ((13'sd3582/*3582:xpc10*/==xpc10))  xpc10 <= 13'sd3583/*3583:xpc10*/;
                  if ((13'sd3583/*3583:xpc10*/==xpc10))  xpc10 <= 13'sd3584/*3584:xpc10*/;
                  if ((13'sd3585/*3585:xpc10*/==xpc10))  xpc10 <= 13'sd698/*698:xpc10*/;
                  if ((13'sd3586/*3586:xpc10*/==xpc10))  xpc10 <= 13'sd3587/*3587:xpc10*/;
                  if ((13'sd3587/*3587:xpc10*/==xpc10))  xpc10 <= 13'sd3588/*3588:xpc10*/;
                  if ((13'sd3590/*3590:xpc10*/==xpc10))  xpc10 <= 13'sd3578/*3578:xpc10*/;
                  if ((13'sd3591/*3591:xpc10*/==xpc10))  xpc10 <= 13'sd3592/*3592:xpc10*/;
                  if ((13'sd3592/*3592:xpc10*/==xpc10))  xpc10 <= 13'sd3593/*3593:xpc10*/;
                  if ((13'sd3594/*3594:xpc10*/==xpc10))  xpc10 <= 13'sd3566/*3566:xpc10*/;
                  if ((13'sd3595/*3595:xpc10*/==xpc10))  xpc10 <= 13'sd3596/*3596:xpc10*/;
                  if ((13'sd3596/*3596:xpc10*/==xpc10))  xpc10 <= 13'sd3597/*3597:xpc10*/;
                  if ((13'sd3598/*3598:xpc10*/==xpc10))  xpc10 <= 13'sd3599/*3599:xpc10*/;
                  if ((13'sd3599/*3599:xpc10*/==xpc10))  xpc10 <= 13'sd3600/*3600:xpc10*/;
                  if ((13'sd3600/*3600:xpc10*/==xpc10))  xpc10 <= 13'sd3601/*3601:xpc10*/;
                  if ((13'sd3601/*3601:xpc10*/==xpc10))  xpc10 <= 13'sd3602/*3602:xpc10*/;
                  if ((13'sd3603/*3603:xpc10*/==xpc10))  xpc10 <= 13'sd3604/*3604:xpc10*/;
                  if ((13'sd3604/*3604:xpc10*/==xpc10))  xpc10 <= 13'sd3605/*3605:xpc10*/;
                  if ((13'sd3605/*3605:xpc10*/==xpc10))  xpc10 <= 13'sd3606/*3606:xpc10*/;
                  if ((13'sd3607/*3607:xpc10*/==xpc10))  xpc10 <= 13'sd3608/*3608:xpc10*/;
                  if ((13'sd3608/*3608:xpc10*/==xpc10))  xpc10 <= 13'sd3609/*3609:xpc10*/;
                  if ((13'sd3609/*3609:xpc10*/==xpc10))  xpc10 <= 13'sd3610/*3610:xpc10*/;
                  if ((13'sd3613/*3613:xpc10*/==xpc10))  xpc10 <= 13'sd3614/*3614:xpc10*/;
                  if ((13'sd3614/*3614:xpc10*/==xpc10))  xpc10 <= 13'sd3615/*3615:xpc10*/;
                  if ((13'sd3615/*3615:xpc10*/==xpc10))  xpc10 <= 13'sd3616/*3616:xpc10*/;
                  if ((13'sd3617/*3617:xpc10*/==xpc10))  xpc10 <= 13'sd3618/*3618:xpc10*/;
                  if ((13'sd3618/*3618:xpc10*/==xpc10))  xpc10 <= 13'sd3619/*3619:xpc10*/;
                  if ((13'sd3619/*3619:xpc10*/==xpc10))  xpc10 <= 13'sd3620/*3620:xpc10*/;
                  if ((13'sd3620/*3620:xpc10*/==xpc10))  xpc10 <= 13'sd3621/*3621:xpc10*/;
                  if ((13'sd3621/*3621:xpc10*/==xpc10))  xpc10 <= 13'sd3622/*3622:xpc10*/;
                  if ((13'sd3622/*3622:xpc10*/==xpc10))  xpc10 <= 13'sd3623/*3623:xpc10*/;
                  if ((13'sd3623/*3623:xpc10*/==xpc10))  xpc10 <= 13'sd3624/*3624:xpc10*/;
                  if ((13'sd3625/*3625:xpc10*/==xpc10))  xpc10 <= 13'sd3626/*3626:xpc10*/;
                  if ((13'sd3626/*3626:xpc10*/==xpc10))  xpc10 <= 13'sd3627/*3627:xpc10*/;
                  if ((13'sd3627/*3627:xpc10*/==xpc10))  xpc10 <= 13'sd3628/*3628:xpc10*/;
                  if ((13'sd3628/*3628:xpc10*/==xpc10))  xpc10 <= 13'sd3629/*3629:xpc10*/;
                  if ((13'sd3629/*3629:xpc10*/==xpc10))  xpc10 <= 13'sd3630/*3630:xpc10*/;
                  if ((13'sd3630/*3630:xpc10*/==xpc10))  xpc10 <= 13'sd3631/*3631:xpc10*/;
                  if ((13'sd3631/*3631:xpc10*/==xpc10))  xpc10 <= 13'sd3632/*3632:xpc10*/;
                  if ((13'sd3634/*3634:xpc10*/==xpc10))  xpc10 <= 13'sd3635/*3635:xpc10*/;
                  if ((13'sd3635/*3635:xpc10*/==xpc10))  xpc10 <= 13'sd3636/*3636:xpc10*/;
                  if ((13'sd3636/*3636:xpc10*/==xpc10))  xpc10 <= 13'sd3637/*3637:xpc10*/;
                  if ((13'sd3638/*3638:xpc10*/==xpc10))  xpc10 <= 13'sd3639/*3639:xpc10*/;
                  if ((13'sd3639/*3639:xpc10*/==xpc10))  xpc10 <= 13'sd3640/*3640:xpc10*/;
                  if ((13'sd3640/*3640:xpc10*/==xpc10))  xpc10 <= 13'sd3641/*3641:xpc10*/;
                  if ((13'sd3642/*3642:xpc10*/==xpc10))  xpc10 <= 13'sd3643/*3643:xpc10*/;
                  if ((13'sd3643/*3643:xpc10*/==xpc10))  xpc10 <= 13'sd3644/*3644:xpc10*/;
                  if ((13'sd3644/*3644:xpc10*/==xpc10))  xpc10 <= 13'sd3645/*3645:xpc10*/;
                  if ((13'sd3646/*3646:xpc10*/==xpc10))  xpc10 <= 13'sd3647/*3647:xpc10*/;
                  if ((13'sd3647/*3647:xpc10*/==xpc10))  xpc10 <= 13'sd3648/*3648:xpc10*/;
                  if ((13'sd3648/*3648:xpc10*/==xpc10))  xpc10 <= 13'sd3649/*3649:xpc10*/;
                  if ((13'sd3650/*3650:xpc10*/==xpc10))  xpc10 <= 13'sd3651/*3651:xpc10*/;
                  if ((13'sd3651/*3651:xpc10*/==xpc10))  xpc10 <= 13'sd3652/*3652:xpc10*/;
                  if ((13'sd3652/*3652:xpc10*/==xpc10))  xpc10 <= 13'sd3653/*3653:xpc10*/;
                  if ((13'sd3654/*3654:xpc10*/==xpc10))  xpc10 <= 13'sd3655/*3655:xpc10*/;
                  if ((13'sd3655/*3655:xpc10*/==xpc10))  xpc10 <= 13'sd3656/*3656:xpc10*/;
                  if ((13'sd3656/*3656:xpc10*/==xpc10))  xpc10 <= 13'sd3657/*3657:xpc10*/;
                  if ((13'sd3658/*3658:xpc10*/==xpc10))  xpc10 <= 13'sd3582/*3582:xpc10*/;
                  if ((13'sd3659/*3659:xpc10*/==xpc10))  xpc10 <= 13'sd3660/*3660:xpc10*/;
                  if ((13'sd3660/*3660:xpc10*/==xpc10))  xpc10 <= 13'sd3661/*3661:xpc10*/;
                  if ((13'sd3662/*3662:xpc10*/==xpc10))  xpc10 <= 13'sd3655/*3655:xpc10*/;
                  if ((13'sd3663/*3663:xpc10*/==xpc10))  xpc10 <= 13'sd3664/*3664:xpc10*/;
                  if ((13'sd3664/*3664:xpc10*/==xpc10))  xpc10 <= 13'sd3665/*3665:xpc10*/;
                  if ((13'sd3666/*3666:xpc10*/==xpc10))  xpc10 <= 13'sd3667/*3667:xpc10*/;
                  if ((13'sd3667/*3667:xpc10*/==xpc10))  xpc10 <= 13'sd3668/*3668:xpc10*/;
                  if ((13'sd3668/*3668:xpc10*/==xpc10))  xpc10 <= 13'sd3669/*3669:xpc10*/;
                  if ((13'sd3673/*3673:xpc10*/==xpc10))  xpc10 <= 13'sd3674/*3674:xpc10*/;
                  if ((13'sd3674/*3674:xpc10*/==xpc10))  xpc10 <= 13'sd3675/*3675:xpc10*/;
                  if ((13'sd3675/*3675:xpc10*/==xpc10))  xpc10 <= 13'sd3676/*3676:xpc10*/;
                  if ((13'sd3678/*3678:xpc10*/==xpc10))  xpc10 <= 13'sd3679/*3679:xpc10*/;
                  if ((13'sd3679/*3679:xpc10*/==xpc10))  xpc10 <= 13'sd3680/*3680:xpc10*/;
                  if ((13'sd3680/*3680:xpc10*/==xpc10))  xpc10 <= 13'sd3681/*3681:xpc10*/;
                  if ((13'sd3682/*3682:xpc10*/==xpc10))  xpc10 <= 13'sd3608/*3608:xpc10*/;
                  if ((13'sd3683/*3683:xpc10*/==xpc10))  xpc10 <= 13'sd3684/*3684:xpc10*/;
                  if ((13'sd3684/*3684:xpc10*/==xpc10))  xpc10 <= 13'sd3685/*3685:xpc10*/;
                  if ((13'sd3687/*3687:xpc10*/==xpc10))  xpc10 <= 13'sd3679/*3679:xpc10*/;
                  if ((13'sd3688/*3688:xpc10*/==xpc10))  xpc10 <= 13'sd3689/*3689:xpc10*/;
                  if ((13'sd3689/*3689:xpc10*/==xpc10))  xpc10 <= 13'sd3690/*3690:xpc10*/;
                  if ((13'sd3691/*3691:xpc10*/==xpc10))  xpc10 <= 13'sd3692/*3692:xpc10*/;
                  if ((13'sd3692/*3692:xpc10*/==xpc10))  xpc10 <= 13'sd3693/*3693:xpc10*/;
                  if ((13'sd3693/*3693:xpc10*/==xpc10))  xpc10 <= 13'sd3694/*3694:xpc10*/;
                  if ((13'sd3695/*3695:xpc10*/==xpc10))  xpc10 <= 13'sd3696/*3696:xpc10*/;
                  if ((13'sd3696/*3696:xpc10*/==xpc10))  xpc10 <= 13'sd3697/*3697:xpc10*/;
                  if ((13'sd3697/*3697:xpc10*/==xpc10))  xpc10 <= 13'sd3698/*3698:xpc10*/;
                  if ((13'sd3699/*3699:xpc10*/==xpc10))  xpc10 <= 13'sd3608/*3608:xpc10*/;
                  if ((13'sd3700/*3700:xpc10*/==xpc10))  xpc10 <= 13'sd3701/*3701:xpc10*/;
                  if ((13'sd3701/*3701:xpc10*/==xpc10))  xpc10 <= 13'sd3702/*3702:xpc10*/;
                  if ((13'sd3703/*3703:xpc10*/==xpc10))  xpc10 <= 13'sd3696/*3696:xpc10*/;
                  if ((13'sd3704/*3704:xpc10*/==xpc10))  xpc10 <= 13'sd3705/*3705:xpc10*/;
                  if ((13'sd3705/*3705:xpc10*/==xpc10))  xpc10 <= 13'sd3706/*3706:xpc10*/;
                  if ((13'sd3708/*3708:xpc10*/==xpc10))  xpc10 <= 13'sd3522/*3522:xpc10*/;
                  if ((13'sd3709/*3709:xpc10*/==xpc10))  xpc10 <= 13'sd3710/*3710:xpc10*/;
                  if ((13'sd3710/*3710:xpc10*/==xpc10))  xpc10 <= 13'sd3711/*3711:xpc10*/;
                  if ((13'sd3713/*3713:xpc10*/==xpc10))  xpc10 <= 13'sd3507/*3507:xpc10*/;
                  if ((13'sd3714/*3714:xpc10*/==xpc10))  xpc10 <= 13'sd3715/*3715:xpc10*/;
                  if ((13'sd3715/*3715:xpc10*/==xpc10))  xpc10 <= 13'sd3716/*3716:xpc10*/;
                  if ((13'sd3718/*3718:xpc10*/==xpc10))  xpc10 <= 13'sd3492/*3492:xpc10*/;
                  if ((13'sd3719/*3719:xpc10*/==xpc10))  xpc10 <= 13'sd3720/*3720:xpc10*/;
                  if ((13'sd3720/*3720:xpc10*/==xpc10))  xpc10 <= 13'sd3721/*3721:xpc10*/;
                  if ((13'sd3721/*3721:xpc10*/==xpc10))  xpc10 <= 13'sd3722/*3722:xpc10*/;
                  if ((13'sd3722/*3722:xpc10*/==xpc10))  xpc10 <= 13'sd3479/*3479:xpc10*/;
                  if ((13'sd3723/*3723:xpc10*/==xpc10))  xpc10 <= 13'sd3724/*3724:xpc10*/;
                  if ((13'sd3724/*3724:xpc10*/==xpc10))  xpc10 <= 13'sd3725/*3725:xpc10*/;
                  if ((13'sd3726/*3726:xpc10*/==xpc10))  xpc10 <= 13'sd3431/*3431:xpc10*/;
                  if ((13'sd3727/*3727:xpc10*/==xpc10))  xpc10 <= 13'sd3728/*3728:xpc10*/;
                  if ((13'sd3728/*3728:xpc10*/==xpc10))  xpc10 <= 13'sd3729/*3729:xpc10*/;
                  if ((13'sd3730/*3730:xpc10*/==xpc10))  xpc10 <= 13'sd3369/*3369:xpc10*/;
                  if ((13'sd3731/*3731:xpc10*/==xpc10))  xpc10 <= 13'sd3732/*3732:xpc10*/;
                  if ((13'sd3732/*3732:xpc10*/==xpc10))  xpc10 <= 13'sd3733/*3733:xpc10*/;
                  if ((13'sd3734/*3734:xpc10*/==xpc10))  xpc10 <= 13'sd637/*637:xpc10*/;
                  if ((13'sd3735/*3735:xpc10*/==xpc10))  xpc10 <= 13'sd3736/*3736:xpc10*/;
                  if ((13'sd3736/*3736:xpc10*/==xpc10))  xpc10 <= 13'sd3737/*3737:xpc10*/;
                  if ((13'sd3738/*3738:xpc10*/==xpc10))  xpc10 <= 13'sd626/*626:xpc10*/;
                  if ((13'sd3739/*3739:xpc10*/==xpc10))  xpc10 <= 13'sd3740/*3740:xpc10*/;
                  if ((13'sd3740/*3740:xpc10*/==xpc10))  xpc10 <= 13'sd3741/*3741:xpc10*/;
                  if ((13'sd3743/*3743:xpc10*/==xpc10))  xpc10 <= 13'sd3744/*3744:xpc10*/;
                  if ((13'sd3744/*3744:xpc10*/==xpc10))  xpc10 <= 13'sd3745/*3745:xpc10*/;
                  if ((13'sd3745/*3745:xpc10*/==xpc10))  xpc10 <= 13'sd3746/*3746:xpc10*/;
                  if ((13'sd3747/*3747:xpc10*/==xpc10))  xpc10 <= 13'sd3748/*3748:xpc10*/;
                  if ((13'sd3748/*3748:xpc10*/==xpc10))  xpc10 <= 13'sd3749/*3749:xpc10*/;
                  if ((13'sd3749/*3749:xpc10*/==xpc10))  xpc10 <= 13'sd3750/*3750:xpc10*/;
                  if ((13'sd3754/*3754:xpc10*/==xpc10))  xpc10 <= 13'sd3755/*3755:xpc10*/;
                  if ((13'sd3755/*3755:xpc10*/==xpc10))  xpc10 <= 13'sd3756/*3756:xpc10*/;
                  if ((13'sd3756/*3756:xpc10*/==xpc10))  xpc10 <= 13'sd3757/*3757:xpc10*/;
                  if ((13'sd3759/*3759:xpc10*/==xpc10))  xpc10 <= 13'sd3760/*3760:xpc10*/;
                  if ((13'sd3760/*3760:xpc10*/==xpc10))  xpc10 <= 13'sd3761/*3761:xpc10*/;
                  if ((13'sd3761/*3761:xpc10*/==xpc10))  xpc10 <= 13'sd3762/*3762:xpc10*/;
                  if ((13'sd3763/*3763:xpc10*/==xpc10))  xpc10 <= 13'sd3764/*3764:xpc10*/;
                  if ((13'sd3764/*3764:xpc10*/==xpc10))  xpc10 <= 13'sd3765/*3765:xpc10*/;
                  if ((13'sd3765/*3765:xpc10*/==xpc10))  xpc10 <= 13'sd3766/*3766:xpc10*/;
                  if ((13'sd3768/*3768:xpc10*/==xpc10))  xpc10 <= 13'sd3769/*3769:xpc10*/;
                  if ((13'sd3769/*3769:xpc10*/==xpc10))  xpc10 <= 13'sd3770/*3770:xpc10*/;
                  if ((13'sd3770/*3770:xpc10*/==xpc10))  xpc10 <= 13'sd3771/*3771:xpc10*/;
                  if ((13'sd3775/*3775:xpc10*/==xpc10))  xpc10 <= 13'sd3776/*3776:xpc10*/;
                  if ((13'sd3776/*3776:xpc10*/==xpc10))  xpc10 <= 13'sd3777/*3777:xpc10*/;
                  if ((13'sd3777/*3777:xpc10*/==xpc10))  xpc10 <= 13'sd3778/*3778:xpc10*/;
                  if ((13'sd3779/*3779:xpc10*/==xpc10))  xpc10 <= 13'sd3780/*3780:xpc10*/;
                  if ((13'sd3780/*3780:xpc10*/==xpc10))  xpc10 <= 13'sd3781/*3781:xpc10*/;
                  if ((13'sd3781/*3781:xpc10*/==xpc10))  xpc10 <= 13'sd3782/*3782:xpc10*/;
                  if ((13'sd3783/*3783:xpc10*/==xpc10))  xpc10 <= 13'sd612/*612:xpc10*/;
                  if ((13'sd3784/*3784:xpc10*/==xpc10))  xpc10 <= 13'sd3785/*3785:xpc10*/;
                  if ((13'sd3785/*3785:xpc10*/==xpc10))  xpc10 <= 13'sd3786/*3786:xpc10*/;
                  if ((13'sd3787/*3787:xpc10*/==xpc10))  xpc10 <= 13'sd3780/*3780:xpc10*/;
                  if ((13'sd3788/*3788:xpc10*/==xpc10))  xpc10 <= 13'sd3789/*3789:xpc10*/;
                  if ((13'sd3789/*3789:xpc10*/==xpc10))  xpc10 <= 13'sd3790/*3790:xpc10*/;
                  if ((13'sd3791/*3791:xpc10*/==xpc10))  xpc10 <= 13'sd3748/*3748:xpc10*/;
                  if ((13'sd3792/*3792:xpc10*/==xpc10))  xpc10 <= 13'sd3793/*3793:xpc10*/;
                  if ((13'sd3793/*3793:xpc10*/==xpc10))  xpc10 <= 13'sd3794/*3794:xpc10*/;
                  if ((13'sd3795/*3795:xpc10*/==xpc10))  xpc10 <= 13'sd3796/*3796:xpc10*/;
                  if ((13'sd3796/*3796:xpc10*/==xpc10))  xpc10 <= 13'sd3797/*3797:xpc10*/;
                  if ((13'sd3797/*3797:xpc10*/==xpc10))  xpc10 <= 13'sd3798/*3798:xpc10*/;
                  if ((13'sd3799/*3799:xpc10*/==xpc10))  xpc10 <= 13'sd600/*600:xpc10*/;
                  if ((13'sd3800/*3800:xpc10*/==xpc10))  xpc10 <= 13'sd3801/*3801:xpc10*/;
                  if ((13'sd3801/*3801:xpc10*/==xpc10))  xpc10 <= 13'sd3802/*3802:xpc10*/;
                  if ((13'sd3803/*3803:xpc10*/==xpc10))  xpc10 <= 13'sd3804/*3804:xpc10*/;
                  if ((13'sd3804/*3804:xpc10*/==xpc10))  xpc10 <= 13'sd3805/*3805:xpc10*/;
                  if ((13'sd3805/*3805:xpc10*/==xpc10))  xpc10 <= 13'sd3806/*3806:xpc10*/;
                  if ((13'sd3807/*3807:xpc10*/==xpc10))  xpc10 <= 13'sd600/*600:xpc10*/;
                  if ((13'sd3808/*3808:xpc10*/==xpc10))  xpc10 <= 13'sd3809/*3809:xpc10*/;
                  if ((13'sd3809/*3809:xpc10*/==xpc10))  xpc10 <= 13'sd3810/*3810:xpc10*/;
                  if ((13'sd3811/*3811:xpc10*/==xpc10))  xpc10 <= 13'sd600/*600:xpc10*/;
                  if ((13'sd3812/*3812:xpc10*/==xpc10))  xpc10 <= 13'sd3813/*3813:xpc10*/;
                  if ((13'sd3813/*3813:xpc10*/==xpc10))  xpc10 <= 13'sd3814/*3814:xpc10*/;
                  if ((13'sd3815/*3815:xpc10*/==xpc10))  xpc10 <= 13'sd581/*581:xpc10*/;
                  if ((13'sd3816/*3816:xpc10*/==xpc10))  xpc10 <= 13'sd3817/*3817:xpc10*/;
                  if ((13'sd3817/*3817:xpc10*/==xpc10))  xpc10 <= 13'sd3818/*3818:xpc10*/;
                  if ((13'sd3819/*3819:xpc10*/==xpc10))  xpc10 <= 13'sd571/*571:xpc10*/;
                  if ((13'sd3820/*3820:xpc10*/==xpc10))  xpc10 <= 13'sd3821/*3821:xpc10*/;
                  if ((13'sd3821/*3821:xpc10*/==xpc10))  xpc10 <= 13'sd3822/*3822:xpc10*/;
                  if ((13'sd3823/*3823:xpc10*/==xpc10))  xpc10 <= 13'sd3824/*3824:xpc10*/;
                  if ((13'sd3824/*3824:xpc10*/==xpc10))  xpc10 <= 13'sd3825/*3825:xpc10*/;
                  if ((13'sd3825/*3825:xpc10*/==xpc10))  xpc10 <= 13'sd3826/*3826:xpc10*/;
                  if ((13'sd3827/*3827:xpc10*/==xpc10))  xpc10 <= 13'sd3828/*3828:xpc10*/;
                  if ((13'sd3828/*3828:xpc10*/==xpc10))  xpc10 <= 13'sd3829/*3829:xpc10*/;
                  if ((13'sd3829/*3829:xpc10*/==xpc10))  xpc10 <= 13'sd3830/*3830:xpc10*/;
                  if ((13'sd3830/*3830:xpc10*/==xpc10))  xpc10 <= 13'sd3831/*3831:xpc10*/;
                  if ((13'sd3832/*3832:xpc10*/==xpc10))  xpc10 <= 13'sd604/*604:xpc10*/;
                  if ((13'sd3833/*3833:xpc10*/==xpc10))  xpc10 <= 13'sd3834/*3834:xpc10*/;
                  if ((13'sd3834/*3834:xpc10*/==xpc10))  xpc10 <= 13'sd3835/*3835:xpc10*/;
                  if ((13'sd3836/*3836:xpc10*/==xpc10))  xpc10 <= 13'sd3837/*3837:xpc10*/;
                  if ((13'sd3837/*3837:xpc10*/==xpc10))  xpc10 <= 13'sd3838/*3838:xpc10*/;
                  if ((13'sd3838/*3838:xpc10*/==xpc10))  xpc10 <= 13'sd3839/*3839:xpc10*/;
                  if ((13'sd3840/*3840:xpc10*/==xpc10))  xpc10 <= 13'sd3841/*3841:xpc10*/;
                  if ((13'sd3841/*3841:xpc10*/==xpc10))  xpc10 <= 13'sd3842/*3842:xpc10*/;
                  if ((13'sd3842/*3842:xpc10*/==xpc10))  xpc10 <= 13'sd3843/*3843:xpc10*/;
                  if ((13'sd3844/*3844:xpc10*/==xpc10))  xpc10 <= 13'sd604/*604:xpc10*/;
                  if ((13'sd3845/*3845:xpc10*/==xpc10))  xpc10 <= 13'sd3846/*3846:xpc10*/;
                  if ((13'sd3846/*3846:xpc10*/==xpc10))  xpc10 <= 13'sd3847/*3847:xpc10*/;
                  if ((13'sd3848/*3848:xpc10*/==xpc10))  xpc10 <= 13'sd3841/*3841:xpc10*/;
                  if ((13'sd3849/*3849:xpc10*/==xpc10))  xpc10 <= 13'sd3850/*3850:xpc10*/;
                  if ((13'sd3850/*3850:xpc10*/==xpc10))  xpc10 <= 13'sd3851/*3851:xpc10*/;
                  if ((13'sd3852/*3852:xpc10*/==xpc10))  xpc10 <= 13'sd3853/*3853:xpc10*/;
                  if ((13'sd3853/*3853:xpc10*/==xpc10))  xpc10 <= 13'sd3854/*3854:xpc10*/;
                  if ((13'sd3854/*3854:xpc10*/==xpc10))  xpc10 <= 13'sd3855/*3855:xpc10*/;
                  if ((13'sd3856/*3856:xpc10*/==xpc10))  xpc10 <= 13'sd3857/*3857:xpc10*/;
                  if ((13'sd3857/*3857:xpc10*/==xpc10))  xpc10 <= 13'sd3858/*3858:xpc10*/;
                  if ((13'sd3858/*3858:xpc10*/==xpc10))  xpc10 <= 13'sd3859/*3859:xpc10*/;
                  if ((13'sd3862/*3862:xpc10*/==xpc10))  xpc10 <= 13'sd3863/*3863:xpc10*/;
                  if ((13'sd3863/*3863:xpc10*/==xpc10))  xpc10 <= 13'sd3864/*3864:xpc10*/;
                  if ((13'sd3864/*3864:xpc10*/==xpc10))  xpc10 <= 13'sd3865/*3865:xpc10*/;
                  if ((13'sd3866/*3866:xpc10*/==xpc10))  xpc10 <= 13'sd3867/*3867:xpc10*/;
                  if ((13'sd3867/*3867:xpc10*/==xpc10))  xpc10 <= 13'sd3868/*3868:xpc10*/;
                  if ((13'sd3868/*3868:xpc10*/==xpc10))  xpc10 <= 13'sd3869/*3869:xpc10*/;
                  if ((13'sd3872/*3872:xpc10*/==xpc10))  xpc10 <= 13'sd3873/*3873:xpc10*/;
                  if ((13'sd3873/*3873:xpc10*/==xpc10))  xpc10 <= 13'sd3874/*3874:xpc10*/;
                  if ((13'sd3874/*3874:xpc10*/==xpc10))  xpc10 <= 13'sd3875/*3875:xpc10*/;
                  if ((13'sd3876/*3876:xpc10*/==xpc10))  xpc10 <= 13'sd3877/*3877:xpc10*/;
                  if ((13'sd3877/*3877:xpc10*/==xpc10))  xpc10 <= 13'sd3878/*3878:xpc10*/;
                  if ((13'sd3878/*3878:xpc10*/==xpc10))  xpc10 <= 13'sd3879/*3879:xpc10*/;
                  if ((13'sd3883/*3883:xpc10*/==xpc10))  xpc10 <= 13'sd3884/*3884:xpc10*/;
                  if ((13'sd3884/*3884:xpc10*/==xpc10))  xpc10 <= 13'sd3885/*3885:xpc10*/;
                  if ((13'sd3885/*3885:xpc10*/==xpc10))  xpc10 <= 13'sd3886/*3886:xpc10*/;
                  if ((13'sd3886/*3886:xpc10*/==xpc10))  xpc10 <= 13'sd3887/*3887:xpc10*/;
                  if ((13'sd3887/*3887:xpc10*/==xpc10))  xpc10 <= 13'sd3888/*3888:xpc10*/;
                  if ((13'sd3888/*3888:xpc10*/==xpc10))  xpc10 <= 13'sd3889/*3889:xpc10*/;
                  if ((13'sd3889/*3889:xpc10*/==xpc10))  xpc10 <= 13'sd3890/*3890:xpc10*/;
                  if ((13'sd3891/*3891:xpc10*/==xpc10))  xpc10 <= 13'sd3892/*3892:xpc10*/;
                  if ((13'sd3892/*3892:xpc10*/==xpc10))  xpc10 <= 13'sd3893/*3893:xpc10*/;
                  if ((13'sd3893/*3893:xpc10*/==xpc10))  xpc10 <= 13'sd3894/*3894:xpc10*/;
                  if ((13'sd3895/*3895:xpc10*/==xpc10))  xpc10 <= 13'sd3896/*3896:xpc10*/;
                  if ((13'sd3896/*3896:xpc10*/==xpc10))  xpc10 <= 13'sd3897/*3897:xpc10*/;
                  if ((13'sd3897/*3897:xpc10*/==xpc10))  xpc10 <= 13'sd3898/*3898:xpc10*/;
                  if ((13'sd3899/*3899:xpc10*/==xpc10))  xpc10 <= 13'sd604/*604:xpc10*/;
                  if ((13'sd3900/*3900:xpc10*/==xpc10))  xpc10 <= 13'sd3901/*3901:xpc10*/;
                  if ((13'sd3901/*3901:xpc10*/==xpc10))  xpc10 <= 13'sd3902/*3902:xpc10*/;
                  if ((13'sd3903/*3903:xpc10*/==xpc10))  xpc10 <= 13'sd3904/*3904:xpc10*/;
                  if ((13'sd3904/*3904:xpc10*/==xpc10))  xpc10 <= 13'sd3905/*3905:xpc10*/;
                  if ((13'sd3905/*3905:xpc10*/==xpc10))  xpc10 <= 13'sd3906/*3906:xpc10*/;
                  if ((13'sd3907/*3907:xpc10*/==xpc10))  xpc10 <= 13'sd3896/*3896:xpc10*/;
                  if ((13'sd3908/*3908:xpc10*/==xpc10))  xpc10 <= 13'sd3909/*3909:xpc10*/;
                  if ((13'sd3909/*3909:xpc10*/==xpc10))  xpc10 <= 13'sd3910/*3910:xpc10*/;
                  if ((13'sd3911/*3911:xpc10*/==xpc10))  xpc10 <= 13'sd3912/*3912:xpc10*/;
                  if ((13'sd3912/*3912:xpc10*/==xpc10))  xpc10 <= 13'sd3913/*3913:xpc10*/;
                  if ((13'sd3913/*3913:xpc10*/==xpc10))  xpc10 <= 13'sd3914/*3914:xpc10*/;
                  if ((13'sd3915/*3915:xpc10*/==xpc10))  xpc10 <= 13'sd3896/*3896:xpc10*/;
                  if ((13'sd3916/*3916:xpc10*/==xpc10))  xpc10 <= 13'sd3917/*3917:xpc10*/;
                  if ((13'sd3917/*3917:xpc10*/==xpc10))  xpc10 <= 13'sd3918/*3918:xpc10*/;
                  if ((13'sd3919/*3919:xpc10*/==xpc10))  xpc10 <= 13'sd3896/*3896:xpc10*/;
                  if ((13'sd3920/*3920:xpc10*/==xpc10))  xpc10 <= 13'sd3921/*3921:xpc10*/;
                  if ((13'sd3921/*3921:xpc10*/==xpc10))  xpc10 <= 13'sd3922/*3922:xpc10*/;
                  if ((13'sd3923/*3923:xpc10*/==xpc10))  xpc10 <= 13'sd3877/*3877:xpc10*/;
                  if ((13'sd3924/*3924:xpc10*/==xpc10))  xpc10 <= 13'sd3925/*3925:xpc10*/;
                  if ((13'sd3925/*3925:xpc10*/==xpc10))  xpc10 <= 13'sd3926/*3926:xpc10*/;
                  if ((13'sd3927/*3927:xpc10*/==xpc10))  xpc10 <= 13'sd3867/*3867:xpc10*/;
                  if ((13'sd3928/*3928:xpc10*/==xpc10))  xpc10 <= 13'sd3929/*3929:xpc10*/;
                  if ((13'sd3929/*3929:xpc10*/==xpc10))  xpc10 <= 13'sd3930/*3930:xpc10*/;
                  if ((13'sd3931/*3931:xpc10*/==xpc10))  xpc10 <= 13'sd3932/*3932:xpc10*/;
                  if ((13'sd3932/*3932:xpc10*/==xpc10))  xpc10 <= 13'sd3933/*3933:xpc10*/;
                  if ((13'sd3933/*3933:xpc10*/==xpc10))  xpc10 <= 13'sd3934/*3934:xpc10*/;
                  if ((13'sd3935/*3935:xpc10*/==xpc10))  xpc10 <= 13'sd3936/*3936:xpc10*/;
                  if ((13'sd3936/*3936:xpc10*/==xpc10))  xpc10 <= 13'sd3937/*3937:xpc10*/;
                  if ((13'sd3937/*3937:xpc10*/==xpc10))  xpc10 <= 13'sd3938/*3938:xpc10*/;
                  if ((13'sd3938/*3938:xpc10*/==xpc10))  xpc10 <= 13'sd3939/*3939:xpc10*/;
                  if ((13'sd3940/*3940:xpc10*/==xpc10))  xpc10 <= 13'sd604/*604:xpc10*/;
                  if ((13'sd3941/*3941:xpc10*/==xpc10))  xpc10 <= 13'sd3942/*3942:xpc10*/;
                  if ((13'sd3942/*3942:xpc10*/==xpc10))  xpc10 <= 13'sd3943/*3943:xpc10*/;
                  if ((13'sd3944/*3944:xpc10*/==xpc10))  xpc10 <= 13'sd3945/*3945:xpc10*/;
                  if ((13'sd3945/*3945:xpc10*/==xpc10))  xpc10 <= 13'sd3946/*3946:xpc10*/;
                  if ((13'sd3946/*3946:xpc10*/==xpc10))  xpc10 <= 13'sd3947/*3947:xpc10*/;
                  if ((13'sd3948/*3948:xpc10*/==xpc10))  xpc10 <= 13'sd3949/*3949:xpc10*/;
                  if ((13'sd3949/*3949:xpc10*/==xpc10))  xpc10 <= 13'sd3950/*3950:xpc10*/;
                  if ((13'sd3950/*3950:xpc10*/==xpc10))  xpc10 <= 13'sd3951/*3951:xpc10*/;
                  if ((13'sd3952/*3952:xpc10*/==xpc10))  xpc10 <= 13'sd604/*604:xpc10*/;
                  if ((13'sd3953/*3953:xpc10*/==xpc10))  xpc10 <= 13'sd3954/*3954:xpc10*/;
                  if ((13'sd3954/*3954:xpc10*/==xpc10))  xpc10 <= 13'sd3955/*3955:xpc10*/;
                  if ((13'sd3956/*3956:xpc10*/==xpc10))  xpc10 <= 13'sd3949/*3949:xpc10*/;
                  if ((13'sd3957/*3957:xpc10*/==xpc10))  xpc10 <= 13'sd3958/*3958:xpc10*/;
                  if ((13'sd3958/*3958:xpc10*/==xpc10))  xpc10 <= 13'sd3959/*3959:xpc10*/;
                  if ((13'sd3960/*3960:xpc10*/==xpc10))  xpc10 <= 13'sd3961/*3961:xpc10*/;
                  if ((13'sd3961/*3961:xpc10*/==xpc10))  xpc10 <= 13'sd3962/*3962:xpc10*/;
                  if ((13'sd3962/*3962:xpc10*/==xpc10))  xpc10 <= 13'sd3963/*3963:xpc10*/;
                  if ((13'sd3964/*3964:xpc10*/==xpc10))  xpc10 <= 13'sd3965/*3965:xpc10*/;
                  if ((13'sd3965/*3965:xpc10*/==xpc10))  xpc10 <= 13'sd3966/*3966:xpc10*/;
                  if ((13'sd3966/*3966:xpc10*/==xpc10))  xpc10 <= 13'sd3967/*3967:xpc10*/;
                  if ((13'sd3968/*3968:xpc10*/==xpc10))  xpc10 <= 13'sd3969/*3969:xpc10*/;
                  if ((13'sd3969/*3969:xpc10*/==xpc10))  xpc10 <= 13'sd3970/*3970:xpc10*/;
                  if ((13'sd3970/*3970:xpc10*/==xpc10))  xpc10 <= 13'sd3971/*3971:xpc10*/;
                  if ((13'sd3972/*3972:xpc10*/==xpc10))  xpc10 <= 13'sd3973/*3973:xpc10*/;
                  if ((13'sd3973/*3973:xpc10*/==xpc10))  xpc10 <= 13'sd3974/*3974:xpc10*/;
                  if ((13'sd3974/*3974:xpc10*/==xpc10))  xpc10 <= 13'sd3975/*3975:xpc10*/;
                  if ((13'sd3976/*3976:xpc10*/==xpc10))  xpc10 <= 13'sd604/*604:xpc10*/;
                  if ((13'sd3977/*3977:xpc10*/==xpc10))  xpc10 <= 13'sd3978/*3978:xpc10*/;
                  if ((13'sd3978/*3978:xpc10*/==xpc10))  xpc10 <= 13'sd3979/*3979:xpc10*/;
                  if ((13'sd3980/*3980:xpc10*/==xpc10))  xpc10 <= 13'sd3973/*3973:xpc10*/;
                  if ((13'sd3981/*3981:xpc10*/==xpc10))  xpc10 <= 13'sd3982/*3982:xpc10*/;
                  if ((13'sd3982/*3982:xpc10*/==xpc10))  xpc10 <= 13'sd3983/*3983:xpc10*/;
                  if ((13'sd3986/*3986:xpc10*/==xpc10))  xpc10 <= 13'sd3987/*3987:xpc10*/;
                  if ((13'sd3987/*3987:xpc10*/==xpc10))  xpc10 <= 13'sd3988/*3988:xpc10*/;
                  if ((13'sd3988/*3988:xpc10*/==xpc10))  xpc10 <= 13'sd3989/*3989:xpc10*/;
                  if ((13'sd3990/*3990:xpc10*/==xpc10))  xpc10 <= 13'sd3991/*3991:xpc10*/;
                  if ((13'sd3991/*3991:xpc10*/==xpc10))  xpc10 <= 13'sd3992/*3992:xpc10*/;
                  if ((13'sd3992/*3992:xpc10*/==xpc10))  xpc10 <= 13'sd3993/*3993:xpc10*/;
                  if ((13'sd3996/*3996:xpc10*/==xpc10))  xpc10 <= 13'sd3997/*3997:xpc10*/;
                  if ((13'sd3997/*3997:xpc10*/==xpc10))  xpc10 <= 13'sd3998/*3998:xpc10*/;
                  if ((13'sd3998/*3998:xpc10*/==xpc10))  xpc10 <= 13'sd3999/*3999:xpc10*/;
                  if ((13'sd4001/*4001:xpc10*/==xpc10))  xpc10 <= 13'sd4002/*4002:xpc10*/;
                  if ((13'sd4002/*4002:xpc10*/==xpc10))  xpc10 <= 13'sd4003/*4003:xpc10*/;
                  if ((13'sd4003/*4003:xpc10*/==xpc10))  xpc10 <= 13'sd4004/*4004:xpc10*/;
                  if ((13'sd4005/*4005:xpc10*/==xpc10))  xpc10 <= 13'sd4006/*4006:xpc10*/;
                  if ((13'sd4006/*4006:xpc10*/==xpc10))  xpc10 <= 13'sd4007/*4007:xpc10*/;
                  if ((13'sd4007/*4007:xpc10*/==xpc10))  xpc10 <= 13'sd4008/*4008:xpc10*/;
                  if ((13'sd4010/*4010:xpc10*/==xpc10))  xpc10 <= 13'sd4011/*4011:xpc10*/;
                  if ((13'sd4011/*4011:xpc10*/==xpc10))  xpc10 <= 13'sd4012/*4012:xpc10*/;
                  if ((13'sd4012/*4012:xpc10*/==xpc10))  xpc10 <= 13'sd4013/*4013:xpc10*/;
                  if ((13'sd4018/*4018:xpc10*/==xpc10))  xpc10 <= 13'sd4019/*4019:xpc10*/;
                  if ((13'sd4019/*4019:xpc10*/==xpc10))  xpc10 <= 13'sd4020/*4020:xpc10*/;
                  if ((13'sd4020/*4020:xpc10*/==xpc10))  xpc10 <= 13'sd4021/*4021:xpc10*/;
                  if ((13'sd4022/*4022:xpc10*/==xpc10))  xpc10 <= 13'sd4023/*4023:xpc10*/;
                  if ((13'sd4023/*4023:xpc10*/==xpc10))  xpc10 <= 13'sd4024/*4024:xpc10*/;
                  if ((13'sd4024/*4024:xpc10*/==xpc10))  xpc10 <= 13'sd4025/*4025:xpc10*/;
                  if ((13'sd4026/*4026:xpc10*/==xpc10))  xpc10 <= 13'sd4027/*4027:xpc10*/;
                  if ((13'sd4027/*4027:xpc10*/==xpc10))  xpc10 <= 13'sd4028/*4028:xpc10*/;
                  if ((13'sd4028/*4028:xpc10*/==xpc10))  xpc10 <= 13'sd4029/*4029:xpc10*/;
                  if ((13'sd4030/*4030:xpc10*/==xpc10))  xpc10 <= 13'sd4031/*4031:xpc10*/;
                  if ((13'sd4031/*4031:xpc10*/==xpc10))  xpc10 <= 13'sd4032/*4032:xpc10*/;
                  if ((13'sd4032/*4032:xpc10*/==xpc10))  xpc10 <= 13'sd4033/*4033:xpc10*/;
                  if ((13'sd4034/*4034:xpc10*/==xpc10))  xpc10 <= 13'sd4035/*4035:xpc10*/;
                  if ((13'sd4035/*4035:xpc10*/==xpc10))  xpc10 <= 13'sd4036/*4036:xpc10*/;
                  if ((13'sd4036/*4036:xpc10*/==xpc10))  xpc10 <= 13'sd4037/*4037:xpc10*/;
                  if ((13'sd4038/*4038:xpc10*/==xpc10))  xpc10 <= 13'sd604/*604:xpc10*/;
                  if ((13'sd4039/*4039:xpc10*/==xpc10))  xpc10 <= 13'sd4040/*4040:xpc10*/;
                  if ((13'sd4040/*4040:xpc10*/==xpc10))  xpc10 <= 13'sd4041/*4041:xpc10*/;
                  if ((13'sd4042/*4042:xpc10*/==xpc10))  xpc10 <= 13'sd4035/*4035:xpc10*/;
                  if ((13'sd4043/*4043:xpc10*/==xpc10))  xpc10 <= 13'sd4044/*4044:xpc10*/;
                  if ((13'sd4044/*4044:xpc10*/==xpc10))  xpc10 <= 13'sd4045/*4045:xpc10*/;
                  if ((13'sd4048/*4048:xpc10*/==xpc10))  xpc10 <= 13'sd4049/*4049:xpc10*/;
                  if ((13'sd4049/*4049:xpc10*/==xpc10))  xpc10 <= 13'sd4050/*4050:xpc10*/;
                  if ((13'sd4050/*4050:xpc10*/==xpc10))  xpc10 <= 13'sd4051/*4051:xpc10*/;
                  if ((13'sd4052/*4052:xpc10*/==xpc10))  xpc10 <= 13'sd4053/*4053:xpc10*/;
                  if ((13'sd4053/*4053:xpc10*/==xpc10))  xpc10 <= 13'sd4054/*4054:xpc10*/;
                  if ((13'sd4054/*4054:xpc10*/==xpc10))  xpc10 <= 13'sd4055/*4055:xpc10*/;
                  if ((13'sd4058/*4058:xpc10*/==xpc10))  xpc10 <= 13'sd4059/*4059:xpc10*/;
                  if ((13'sd4059/*4059:xpc10*/==xpc10))  xpc10 <= 13'sd4060/*4060:xpc10*/;
                  if ((13'sd4060/*4060:xpc10*/==xpc10))  xpc10 <= 13'sd4061/*4061:xpc10*/;
                  if ((13'sd4063/*4063:xpc10*/==xpc10))  xpc10 <= 13'sd4064/*4064:xpc10*/;
                  if ((13'sd4064/*4064:xpc10*/==xpc10))  xpc10 <= 13'sd4065/*4065:xpc10*/;
                  if ((13'sd4065/*4065:xpc10*/==xpc10))  xpc10 <= 13'sd4066/*4066:xpc10*/;
                  if ((13'sd4067/*4067:xpc10*/==xpc10))  xpc10 <= 13'sd4068/*4068:xpc10*/;
                  if ((13'sd4068/*4068:xpc10*/==xpc10))  xpc10 <= 13'sd4069/*4069:xpc10*/;
                  if ((13'sd4069/*4069:xpc10*/==xpc10))  xpc10 <= 13'sd4070/*4070:xpc10*/;
                  if ((13'sd4072/*4072:xpc10*/==xpc10))  xpc10 <= 13'sd4073/*4073:xpc10*/;
                  if ((13'sd4073/*4073:xpc10*/==xpc10))  xpc10 <= 13'sd4074/*4074:xpc10*/;
                  if ((13'sd4074/*4074:xpc10*/==xpc10))  xpc10 <= 13'sd4075/*4075:xpc10*/;
                  if ((13'sd4080/*4080:xpc10*/==xpc10))  xpc10 <= 13'sd4081/*4081:xpc10*/;
                  if ((13'sd4081/*4081:xpc10*/==xpc10))  xpc10 <= 13'sd4082/*4082:xpc10*/;
                  if ((13'sd4082/*4082:xpc10*/==xpc10))  xpc10 <= 13'sd4083/*4083:xpc10*/;
                  if ((13'sd4096/*4096:xpc10*/==xpc10))  xpc10 <= 13'sd4097/*4097:xpc10*/;
                  if ((13'sd4097/*4097:xpc10*/==xpc10))  xpc10 <= 13'sd4098/*4098:xpc10*/;
                  if ((13'sd4098/*4098:xpc10*/==xpc10))  xpc10 <= 13'sd4099/*4099:xpc10*/;
                  if ((13'sd4099/*4099:xpc10*/==xpc10))  xpc10 <= 13'sd4100/*4100:xpc10*/;
                  if ((13'sd4100/*4100:xpc10*/==xpc10))  xpc10 <= 13'sd4101/*4101:xpc10*/;
                  if ((13'sd4101/*4101:xpc10*/==xpc10))  xpc10 <= 13'sd4102/*4102:xpc10*/;
                  if ((13'sd4102/*4102:xpc10*/==xpc10))  xpc10 <= 13'sd4103/*4103:xpc10*/;
                  if ((13'sd4103/*4103:xpc10*/==xpc10))  xpc10 <= 13'sd4104/*4104:xpc10*/;
                  if ((13'sd4108/*4108:xpc10*/==xpc10))  xpc10 <= 13'sd4109/*4109:xpc10*/;
                  if ((13'sd4109/*4109:xpc10*/==xpc10))  xpc10 <= 13'sd4110/*4110:xpc10*/;
                  if ((13'sd4110/*4110:xpc10*/==xpc10))  xpc10 <= 13'sd4111/*4111:xpc10*/;
                  if ((13'sd4113/*4113:xpc10*/==xpc10))  xpc10 <= 13'sd4114/*4114:xpc10*/;
                  if ((13'sd4114/*4114:xpc10*/==xpc10))  xpc10 <= 13'sd4115/*4115:xpc10*/;
                  if ((13'sd4115/*4115:xpc10*/==xpc10))  xpc10 <= 13'sd4116/*4116:xpc10*/;
                  if ((13'sd4123/*4123:xpc10*/==xpc10))  xpc10 <= 13'sd4124/*4124:xpc10*/;
                  if ((13'sd4124/*4124:xpc10*/==xpc10))  xpc10 <= 13'sd4125/*4125:xpc10*/;
                  if ((13'sd4125/*4125:xpc10*/==xpc10))  xpc10 <= 13'sd4126/*4126:xpc10*/;
                  if ((13'sd4128/*4128:xpc10*/==xpc10))  xpc10 <= 13'sd4129/*4129:xpc10*/;
                  if ((13'sd4129/*4129:xpc10*/==xpc10))  xpc10 <= 13'sd4130/*4130:xpc10*/;
                  if ((13'sd4130/*4130:xpc10*/==xpc10))  xpc10 <= 13'sd4131/*4131:xpc10*/;
                  if ((13'sd4138/*4138:xpc10*/==xpc10))  xpc10 <= 13'sd4139/*4139:xpc10*/;
                  if ((13'sd4139/*4139:xpc10*/==xpc10))  xpc10 <= 13'sd4140/*4140:xpc10*/;
                  if ((13'sd4140/*4140:xpc10*/==xpc10))  xpc10 <= 13'sd4141/*4141:xpc10*/;
                  if ((13'sd4143/*4143:xpc10*/==xpc10))  xpc10 <= 13'sd4144/*4144:xpc10*/;
                  if ((13'sd4144/*4144:xpc10*/==xpc10))  xpc10 <= 13'sd4145/*4145:xpc10*/;
                  if ((13'sd4145/*4145:xpc10*/==xpc10))  xpc10 <= 13'sd4146/*4146:xpc10*/;
                  if ((13'sd4148/*4148:xpc10*/==xpc10))  xpc10 <= 13'sd4149/*4149:xpc10*/;
                  if ((13'sd4149/*4149:xpc10*/==xpc10))  xpc10 <= 13'sd4150/*4150:xpc10*/;
                  if ((13'sd4150/*4150:xpc10*/==xpc10))  xpc10 <= 13'sd4151/*4151:xpc10*/;
                  if ((13'sd4153/*4153:xpc10*/==xpc10))  xpc10 <= 13'sd4154/*4154:xpc10*/;
                  if ((13'sd4154/*4154:xpc10*/==xpc10))  xpc10 <= 13'sd4155/*4155:xpc10*/;
                  if ((13'sd4155/*4155:xpc10*/==xpc10))  xpc10 <= 13'sd4156/*4156:xpc10*/;
                  if ((13'sd4158/*4158:xpc10*/==xpc10))  xpc10 <= 13'sd4159/*4159:xpc10*/;
                  if ((13'sd4159/*4159:xpc10*/==xpc10))  xpc10 <= 13'sd4160/*4160:xpc10*/;
                  if ((13'sd4161/*4161:xpc10*/==xpc10))  xpc10 <= 13'sd4162/*4162:xpc10*/;
                  if ((13'sd4162/*4162:xpc10*/==xpc10))  xpc10 <= 13'sd4163/*4163:xpc10*/;
                  if ((13'sd4163/*4163:xpc10*/==xpc10))  xpc10 <= 13'sd4164/*4164:xpc10*/;
                  if ((13'sd4166/*4166:xpc10*/==xpc10))  xpc10 <= 13'sd4167/*4167:xpc10*/;
                  if ((13'sd4167/*4167:xpc10*/==xpc10))  xpc10 <= 13'sd4168/*4168:xpc10*/;
                  if ((13'sd4168/*4168:xpc10*/==xpc10))  xpc10 <= 13'sd4169/*4169:xpc10*/;
                  if ((13'sd4170/*4170:xpc10*/==xpc10))  xpc10 <= 13'sd4171/*4171:xpc10*/;
                  if ((13'sd4171/*4171:xpc10*/==xpc10))  xpc10 <= 13'sd4172/*4172:xpc10*/;
                  if ((13'sd4172/*4172:xpc10*/==xpc10))  xpc10 <= 13'sd4173/*4173:xpc10*/;
                  if ((13'sd4174/*4174:xpc10*/==xpc10))  xpc10 <= 13'sd4175/*4175:xpc10*/;
                  if ((13'sd4175/*4175:xpc10*/==xpc10))  xpc10 <= 13'sd4176/*4176:xpc10*/;
                  if ((13'sd4176/*4176:xpc10*/==xpc10))  xpc10 <= 13'sd4177/*4177:xpc10*/;
                  if ((13'sd4178/*4178:xpc10*/==xpc10))  xpc10 <= 13'sd4179/*4179:xpc10*/;
                  if ((13'sd4179/*4179:xpc10*/==xpc10))  xpc10 <= 13'sd4180/*4180:xpc10*/;
                  if ((13'sd4180/*4180:xpc10*/==xpc10))  xpc10 <= 13'sd4181/*4181:xpc10*/;
                  if ((13'sd4181/*4181:xpc10*/==xpc10))  xpc10 <= 13'sd4182/*4182:xpc10*/;
                  if ((13'sd4183/*4183:xpc10*/==xpc10))  xpc10 <= 13'sd4184/*4184:xpc10*/;
                  if ((13'sd4184/*4184:xpc10*/==xpc10))  xpc10 <= 13'sd4185/*4185:xpc10*/;
                  if ((13'sd4185/*4185:xpc10*/==xpc10))  xpc10 <= 13'sd4186/*4186:xpc10*/;
                  if ((13'sd4187/*4187:xpc10*/==xpc10))  xpc10 <= 13'sd4188/*4188:xpc10*/;
                  if ((13'sd4188/*4188:xpc10*/==xpc10))  xpc10 <= 13'sd4189/*4189:xpc10*/;
                  if ((13'sd4189/*4189:xpc10*/==xpc10))  xpc10 <= 13'sd4190/*4190:xpc10*/;
                  if ((13'sd4194/*4194:xpc10*/==xpc10))  xpc10 <= 13'sd4195/*4195:xpc10*/;
                  if ((13'sd4195/*4195:xpc10*/==xpc10))  xpc10 <= 13'sd4196/*4196:xpc10*/;
                  if ((13'sd4196/*4196:xpc10*/==xpc10))  xpc10 <= 13'sd4197/*4197:xpc10*/;
                  if ((13'sd4199/*4199:xpc10*/==xpc10))  xpc10 <= 13'sd4200/*4200:xpc10*/;
                  if ((13'sd4200/*4200:xpc10*/==xpc10))  xpc10 <= 13'sd4201/*4201:xpc10*/;
                  if ((13'sd4201/*4201:xpc10*/==xpc10))  xpc10 <= 13'sd4202/*4202:xpc10*/;
                  if ((13'sd4203/*4203:xpc10*/==xpc10))  xpc10 <= 13'sd4204/*4204:xpc10*/;
                  if ((13'sd4204/*4204:xpc10*/==xpc10))  xpc10 <= 13'sd4205/*4205:xpc10*/;
                  if ((13'sd4205/*4205:xpc10*/==xpc10))  xpc10 <= 13'sd4206/*4206:xpc10*/;
                  if ((13'sd4207/*4207:xpc10*/==xpc10))  xpc10 <= 13'sd604/*604:xpc10*/;
                  if ((13'sd4208/*4208:xpc10*/==xpc10))  xpc10 <= 13'sd4209/*4209:xpc10*/;
                  if ((13'sd4209/*4209:xpc10*/==xpc10))  xpc10 <= 13'sd4210/*4210:xpc10*/;
                  if ((13'sd4212/*4212:xpc10*/==xpc10))  xpc10 <= 13'sd4200/*4200:xpc10*/;
                  if ((13'sd4213/*4213:xpc10*/==xpc10))  xpc10 <= 13'sd4214/*4214:xpc10*/;
                  if ((13'sd4214/*4214:xpc10*/==xpc10))  xpc10 <= 13'sd4215/*4215:xpc10*/;
                  if ((13'sd4216/*4216:xpc10*/==xpc10))  xpc10 <= 13'sd4188/*4188:xpc10*/;
                  if ((13'sd4217/*4217:xpc10*/==xpc10))  xpc10 <= 13'sd4218/*4218:xpc10*/;
                  if ((13'sd4218/*4218:xpc10*/==xpc10))  xpc10 <= 13'sd4219/*4219:xpc10*/;
                  if ((13'sd4220/*4220:xpc10*/==xpc10))  xpc10 <= 13'sd4221/*4221:xpc10*/;
                  if ((13'sd4221/*4221:xpc10*/==xpc10))  xpc10 <= 13'sd4222/*4222:xpc10*/;
                  if ((13'sd4222/*4222:xpc10*/==xpc10))  xpc10 <= 13'sd4223/*4223:xpc10*/;
                  if ((13'sd4223/*4223:xpc10*/==xpc10))  xpc10 <= 13'sd4224/*4224:xpc10*/;
                  if ((13'sd4225/*4225:xpc10*/==xpc10))  xpc10 <= 13'sd4226/*4226:xpc10*/;
                  if ((13'sd4226/*4226:xpc10*/==xpc10))  xpc10 <= 13'sd4227/*4227:xpc10*/;
                  if ((13'sd4227/*4227:xpc10*/==xpc10))  xpc10 <= 13'sd4228/*4228:xpc10*/;
                  if ((13'sd4229/*4229:xpc10*/==xpc10))  xpc10 <= 13'sd4230/*4230:xpc10*/;
                  if ((13'sd4230/*4230:xpc10*/==xpc10))  xpc10 <= 13'sd4231/*4231:xpc10*/;
                  if ((13'sd4231/*4231:xpc10*/==xpc10))  xpc10 <= 13'sd4232/*4232:xpc10*/;
                  if ((13'sd4235/*4235:xpc10*/==xpc10))  xpc10 <= 13'sd4236/*4236:xpc10*/;
                  if ((13'sd4236/*4236:xpc10*/==xpc10))  xpc10 <= 13'sd4237/*4237:xpc10*/;
                  if ((13'sd4237/*4237:xpc10*/==xpc10))  xpc10 <= 13'sd4238/*4238:xpc10*/;
                  if ((13'sd4239/*4239:xpc10*/==xpc10))  xpc10 <= 13'sd4240/*4240:xpc10*/;
                  if ((13'sd4240/*4240:xpc10*/==xpc10))  xpc10 <= 13'sd4241/*4241:xpc10*/;
                  if ((13'sd4241/*4241:xpc10*/==xpc10))  xpc10 <= 13'sd4242/*4242:xpc10*/;
                  if ((13'sd4242/*4242:xpc10*/==xpc10))  xpc10 <= 13'sd4243/*4243:xpc10*/;
                  if ((13'sd4243/*4243:xpc10*/==xpc10))  xpc10 <= 13'sd4244/*4244:xpc10*/;
                  if ((13'sd4244/*4244:xpc10*/==xpc10))  xpc10 <= 13'sd4245/*4245:xpc10*/;
                  if ((13'sd4245/*4245:xpc10*/==xpc10))  xpc10 <= 13'sd4246/*4246:xpc10*/;
                  if ((13'sd4247/*4247:xpc10*/==xpc10))  xpc10 <= 13'sd4248/*4248:xpc10*/;
                  if ((13'sd4248/*4248:xpc10*/==xpc10))  xpc10 <= 13'sd4249/*4249:xpc10*/;
                  if ((13'sd4249/*4249:xpc10*/==xpc10))  xpc10 <= 13'sd4250/*4250:xpc10*/;
                  if ((13'sd4250/*4250:xpc10*/==xpc10))  xpc10 <= 13'sd4251/*4251:xpc10*/;
                  if ((13'sd4251/*4251:xpc10*/==xpc10))  xpc10 <= 13'sd4252/*4252:xpc10*/;
                  if ((13'sd4252/*4252:xpc10*/==xpc10))  xpc10 <= 13'sd4253/*4253:xpc10*/;
                  if ((13'sd4253/*4253:xpc10*/==xpc10))  xpc10 <= 13'sd4254/*4254:xpc10*/;
                  if ((13'sd4256/*4256:xpc10*/==xpc10))  xpc10 <= 13'sd4257/*4257:xpc10*/;
                  if ((13'sd4257/*4257:xpc10*/==xpc10))  xpc10 <= 13'sd4258/*4258:xpc10*/;
                  if ((13'sd4258/*4258:xpc10*/==xpc10))  xpc10 <= 13'sd4259/*4259:xpc10*/;
                  if ((13'sd4260/*4260:xpc10*/==xpc10))  xpc10 <= 13'sd4261/*4261:xpc10*/;
                  if ((13'sd4261/*4261:xpc10*/==xpc10))  xpc10 <= 13'sd4262/*4262:xpc10*/;
                  if ((13'sd4262/*4262:xpc10*/==xpc10))  xpc10 <= 13'sd4263/*4263:xpc10*/;
                  if ((13'sd4264/*4264:xpc10*/==xpc10))  xpc10 <= 13'sd4265/*4265:xpc10*/;
                  if ((13'sd4265/*4265:xpc10*/==xpc10))  xpc10 <= 13'sd4266/*4266:xpc10*/;
                  if ((13'sd4266/*4266:xpc10*/==xpc10))  xpc10 <= 13'sd4267/*4267:xpc10*/;
                  if ((13'sd4268/*4268:xpc10*/==xpc10))  xpc10 <= 13'sd4269/*4269:xpc10*/;
                  if ((13'sd4269/*4269:xpc10*/==xpc10))  xpc10 <= 13'sd4270/*4270:xpc10*/;
                  if ((13'sd4270/*4270:xpc10*/==xpc10))  xpc10 <= 13'sd4271/*4271:xpc10*/;
                  if ((13'sd4272/*4272:xpc10*/==xpc10))  xpc10 <= 13'sd4273/*4273:xpc10*/;
                  if ((13'sd4273/*4273:xpc10*/==xpc10))  xpc10 <= 13'sd4274/*4274:xpc10*/;
                  if ((13'sd4274/*4274:xpc10*/==xpc10))  xpc10 <= 13'sd4275/*4275:xpc10*/;
                  if ((13'sd4276/*4276:xpc10*/==xpc10))  xpc10 <= 13'sd4277/*4277:xpc10*/;
                  if ((13'sd4277/*4277:xpc10*/==xpc10))  xpc10 <= 13'sd4278/*4278:xpc10*/;
                  if ((13'sd4278/*4278:xpc10*/==xpc10))  xpc10 <= 13'sd4279/*4279:xpc10*/;
                  if ((13'sd4280/*4280:xpc10*/==xpc10))  xpc10 <= 13'sd4204/*4204:xpc10*/;
                  if ((13'sd4281/*4281:xpc10*/==xpc10))  xpc10 <= 13'sd4282/*4282:xpc10*/;
                  if ((13'sd4282/*4282:xpc10*/==xpc10))  xpc10 <= 13'sd4283/*4283:xpc10*/;
                  if ((13'sd4284/*4284:xpc10*/==xpc10))  xpc10 <= 13'sd4277/*4277:xpc10*/;
                  if ((13'sd4285/*4285:xpc10*/==xpc10))  xpc10 <= 13'sd4286/*4286:xpc10*/;
                  if ((13'sd4286/*4286:xpc10*/==xpc10))  xpc10 <= 13'sd4287/*4287:xpc10*/;
                  if ((13'sd4288/*4288:xpc10*/==xpc10))  xpc10 <= 13'sd4289/*4289:xpc10*/;
                  if ((13'sd4289/*4289:xpc10*/==xpc10))  xpc10 <= 13'sd4290/*4290:xpc10*/;
                  if ((13'sd4290/*4290:xpc10*/==xpc10))  xpc10 <= 13'sd4291/*4291:xpc10*/;
                  if ((13'sd4295/*4295:xpc10*/==xpc10))  xpc10 <= 13'sd4296/*4296:xpc10*/;
                  if ((13'sd4296/*4296:xpc10*/==xpc10))  xpc10 <= 13'sd4297/*4297:xpc10*/;
                  if ((13'sd4297/*4297:xpc10*/==xpc10))  xpc10 <= 13'sd4298/*4298:xpc10*/;
                  if ((13'sd4300/*4300:xpc10*/==xpc10))  xpc10 <= 13'sd4301/*4301:xpc10*/;
                  if ((13'sd4301/*4301:xpc10*/==xpc10))  xpc10 <= 13'sd4302/*4302:xpc10*/;
                  if ((13'sd4302/*4302:xpc10*/==xpc10))  xpc10 <= 13'sd4303/*4303:xpc10*/;
                  if ((13'sd4304/*4304:xpc10*/==xpc10))  xpc10 <= 13'sd4230/*4230:xpc10*/;
                  if ((13'sd4305/*4305:xpc10*/==xpc10))  xpc10 <= 13'sd4306/*4306:xpc10*/;
                  if ((13'sd4306/*4306:xpc10*/==xpc10))  xpc10 <= 13'sd4307/*4307:xpc10*/;
                  if ((13'sd4309/*4309:xpc10*/==xpc10))  xpc10 <= 13'sd4301/*4301:xpc10*/;
                  if ((13'sd4310/*4310:xpc10*/==xpc10))  xpc10 <= 13'sd4311/*4311:xpc10*/;
                  if ((13'sd4311/*4311:xpc10*/==xpc10))  xpc10 <= 13'sd4312/*4312:xpc10*/;
                  if ((13'sd4313/*4313:xpc10*/==xpc10))  xpc10 <= 13'sd4314/*4314:xpc10*/;
                  if ((13'sd4314/*4314:xpc10*/==xpc10))  xpc10 <= 13'sd4315/*4315:xpc10*/;
                  if ((13'sd4315/*4315:xpc10*/==xpc10))  xpc10 <= 13'sd4316/*4316:xpc10*/;
                  if ((13'sd4317/*4317:xpc10*/==xpc10))  xpc10 <= 13'sd4318/*4318:xpc10*/;
                  if ((13'sd4318/*4318:xpc10*/==xpc10))  xpc10 <= 13'sd4319/*4319:xpc10*/;
                  if ((13'sd4319/*4319:xpc10*/==xpc10))  xpc10 <= 13'sd4320/*4320:xpc10*/;
                  if ((13'sd4321/*4321:xpc10*/==xpc10))  xpc10 <= 13'sd4230/*4230:xpc10*/;
                  if ((13'sd4322/*4322:xpc10*/==xpc10))  xpc10 <= 13'sd4323/*4323:xpc10*/;
                  if ((13'sd4323/*4323:xpc10*/==xpc10))  xpc10 <= 13'sd4324/*4324:xpc10*/;
                  if ((13'sd4325/*4325:xpc10*/==xpc10))  xpc10 <= 13'sd4318/*4318:xpc10*/;
                  if ((13'sd4326/*4326:xpc10*/==xpc10))  xpc10 <= 13'sd4327/*4327:xpc10*/;
                  if ((13'sd4327/*4327:xpc10*/==xpc10))  xpc10 <= 13'sd4328/*4328:xpc10*/;
                  if ((13'sd4330/*4330:xpc10*/==xpc10))  xpc10 <= 13'sd4144/*4144:xpc10*/;
                  if ((13'sd4331/*4331:xpc10*/==xpc10))  xpc10 <= 13'sd4332/*4332:xpc10*/;
                  if ((13'sd4332/*4332:xpc10*/==xpc10))  xpc10 <= 13'sd4333/*4333:xpc10*/;
                  if ((13'sd4335/*4335:xpc10*/==xpc10))  xpc10 <= 13'sd4129/*4129:xpc10*/;
                  if ((13'sd4336/*4336:xpc10*/==xpc10))  xpc10 <= 13'sd4337/*4337:xpc10*/;
                  if ((13'sd4337/*4337:xpc10*/==xpc10))  xpc10 <= 13'sd4338/*4338:xpc10*/;
                  if ((13'sd4340/*4340:xpc10*/==xpc10))  xpc10 <= 13'sd4114/*4114:xpc10*/;
                  if ((13'sd4341/*4341:xpc10*/==xpc10))  xpc10 <= 13'sd4342/*4342:xpc10*/;
                  if ((13'sd4342/*4342:xpc10*/==xpc10))  xpc10 <= 13'sd4343/*4343:xpc10*/;
                  if ((13'sd4343/*4343:xpc10*/==xpc10))  xpc10 <= 13'sd4344/*4344:xpc10*/;
                  if ((13'sd4344/*4344:xpc10*/==xpc10))  xpc10 <= 13'sd4101/*4101:xpc10*/;
                  if ((13'sd4345/*4345:xpc10*/==xpc10))  xpc10 <= 13'sd4346/*4346:xpc10*/;
                  if ((13'sd4346/*4346:xpc10*/==xpc10))  xpc10 <= 13'sd4347/*4347:xpc10*/;
                  if ((13'sd4348/*4348:xpc10*/==xpc10))  xpc10 <= 13'sd4053/*4053:xpc10*/;
                  if ((13'sd4349/*4349:xpc10*/==xpc10))  xpc10 <= 13'sd4350/*4350:xpc10*/;
                  if ((13'sd4350/*4350:xpc10*/==xpc10))  xpc10 <= 13'sd4351/*4351:xpc10*/;
                  if ((13'sd4352/*4352:xpc10*/==xpc10))  xpc10 <= 13'sd3991/*3991:xpc10*/;
                  if ((13'sd4353/*4353:xpc10*/==xpc10))  xpc10 <= 13'sd4354/*4354:xpc10*/;
                  if ((13'sd4354/*4354:xpc10*/==xpc10))  xpc10 <= 13'sd4355/*4355:xpc10*/;
                  if ((13'sd4356/*4356:xpc10*/==xpc10))  xpc10 <= 13'sd543/*543:xpc10*/;
                  if ((13'sd4357/*4357:xpc10*/==xpc10))  xpc10 <= 13'sd4358/*4358:xpc10*/;
                  if ((13'sd4358/*4358:xpc10*/==xpc10))  xpc10 <= 13'sd4359/*4359:xpc10*/;
                  if ((13'sd4360/*4360:xpc10*/==xpc10))  xpc10 <= 13'sd532/*532:xpc10*/;
                  if ((13'sd4361/*4361:xpc10*/==xpc10))  xpc10 <= 13'sd4362/*4362:xpc10*/;
                  if ((13'sd4362/*4362:xpc10*/==xpc10))  xpc10 <= 13'sd4363/*4363:xpc10*/;
                  if ((13'sd4364/*4364:xpc10*/==xpc10))  xpc10 <= 13'sd4365/*4365:xpc10*/;
                  if ((13'sd4365/*4365:xpc10*/==xpc10))  xpc10 <= 13'sd4366/*4366:xpc10*/;
                  if ((13'sd4366/*4366:xpc10*/==xpc10))  xpc10 <= 13'sd4367/*4367:xpc10*/;
                  if ((13'sd4368/*4368:xpc10*/==xpc10))  xpc10 <= 13'sd507/*507:xpc10*/;
                  if ((13'sd4369/*4369:xpc10*/==xpc10))  xpc10 <= 13'sd4370/*4370:xpc10*/;
                  if ((13'sd4370/*4370:xpc10*/==xpc10))  xpc10 <= 13'sd4371/*4371:xpc10*/;
                  if ((13'sd4372/*4372:xpc10*/==xpc10))  xpc10 <= 13'sd4373/*4373:xpc10*/;
                  if ((13'sd4373/*4373:xpc10*/==xpc10))  xpc10 <= 13'sd4374/*4374:xpc10*/;
                  if ((13'sd4374/*4374:xpc10*/==xpc10))  xpc10 <= 13'sd4375/*4375:xpc10*/;
                  if ((13'sd4376/*4376:xpc10*/==xpc10))  xpc10 <= 13'sd507/*507:xpc10*/;
                  if ((13'sd4377/*4377:xpc10*/==xpc10))  xpc10 <= 13'sd4378/*4378:xpc10*/;
                  if ((13'sd4378/*4378:xpc10*/==xpc10))  xpc10 <= 13'sd4379/*4379:xpc10*/;
                  if ((13'sd4380/*4380:xpc10*/==xpc10))  xpc10 <= 13'sd507/*507:xpc10*/;
                  if ((13'sd4381/*4381:xpc10*/==xpc10))  xpc10 <= 13'sd4382/*4382:xpc10*/;
                  if ((13'sd4382/*4382:xpc10*/==xpc10))  xpc10 <= 13'sd4383/*4383:xpc10*/;
                  if ((13'sd4384/*4384:xpc10*/==xpc10))  xpc10 <= 13'sd488/*488:xpc10*/;
                  if ((13'sd4385/*4385:xpc10*/==xpc10))  xpc10 <= 13'sd4386/*4386:xpc10*/;
                  if ((13'sd4386/*4386:xpc10*/==xpc10))  xpc10 <= 13'sd4387/*4387:xpc10*/;
                  if ((13'sd4388/*4388:xpc10*/==xpc10))  xpc10 <= 13'sd478/*478:xpc10*/;
                  if ((13'sd4389/*4389:xpc10*/==xpc10))  xpc10 <= 13'sd4390/*4390:xpc10*/;
                  if ((13'sd4390/*4390:xpc10*/==xpc10))  xpc10 <= 13'sd4391/*4391:xpc10*/;
                  if ((13'sd4392/*4392:xpc10*/==xpc10))  xpc10 <= 13'sd4393/*4393:xpc10*/;
                  if ((13'sd4393/*4393:xpc10*/==xpc10))  xpc10 <= 13'sd4394/*4394:xpc10*/;
                  if ((13'sd4394/*4394:xpc10*/==xpc10))  xpc10 <= 13'sd4395/*4395:xpc10*/;
                  if ((13'sd4396/*4396:xpc10*/==xpc10))  xpc10 <= 13'sd4397/*4397:xpc10*/;
                  if ((13'sd4397/*4397:xpc10*/==xpc10))  xpc10 <= 13'sd4398/*4398:xpc10*/;
                  if ((13'sd4398/*4398:xpc10*/==xpc10))  xpc10 <= 13'sd4399/*4399:xpc10*/;
                  if ((13'sd4399/*4399:xpc10*/==xpc10))  xpc10 <= 13'sd4400/*4400:xpc10*/;
                  if ((13'sd4401/*4401:xpc10*/==xpc10))  xpc10 <= 13'sd511/*511:xpc10*/;
                  if ((13'sd4402/*4402:xpc10*/==xpc10))  xpc10 <= 13'sd4403/*4403:xpc10*/;
                  if ((13'sd4403/*4403:xpc10*/==xpc10))  xpc10 <= 13'sd4404/*4404:xpc10*/;
                  if ((13'sd4405/*4405:xpc10*/==xpc10))  xpc10 <= 13'sd4406/*4406:xpc10*/;
                  if ((13'sd4406/*4406:xpc10*/==xpc10))  xpc10 <= 13'sd4407/*4407:xpc10*/;
                  if ((13'sd4407/*4407:xpc10*/==xpc10))  xpc10 <= 13'sd4408/*4408:xpc10*/;
                  if ((13'sd4409/*4409:xpc10*/==xpc10))  xpc10 <= 13'sd4410/*4410:xpc10*/;
                  if ((13'sd4410/*4410:xpc10*/==xpc10))  xpc10 <= 13'sd4411/*4411:xpc10*/;
                  if ((13'sd4411/*4411:xpc10*/==xpc10))  xpc10 <= 13'sd4412/*4412:xpc10*/;
                  if ((13'sd4413/*4413:xpc10*/==xpc10))  xpc10 <= 13'sd511/*511:xpc10*/;
                  if ((13'sd4414/*4414:xpc10*/==xpc10))  xpc10 <= 13'sd4415/*4415:xpc10*/;
                  if ((13'sd4415/*4415:xpc10*/==xpc10))  xpc10 <= 13'sd4416/*4416:xpc10*/;
                  if ((13'sd4417/*4417:xpc10*/==xpc10))  xpc10 <= 13'sd4410/*4410:xpc10*/;
                  if ((13'sd4418/*4418:xpc10*/==xpc10))  xpc10 <= 13'sd4419/*4419:xpc10*/;
                  if ((13'sd4419/*4419:xpc10*/==xpc10))  xpc10 <= 13'sd4420/*4420:xpc10*/;
                  if ((13'sd4421/*4421:xpc10*/==xpc10))  xpc10 <= 13'sd4422/*4422:xpc10*/;
                  if ((13'sd4422/*4422:xpc10*/==xpc10))  xpc10 <= 13'sd4423/*4423:xpc10*/;
                  if ((13'sd4423/*4423:xpc10*/==xpc10))  xpc10 <= 13'sd4424/*4424:xpc10*/;
                  if ((13'sd4425/*4425:xpc10*/==xpc10))  xpc10 <= 13'sd4426/*4426:xpc10*/;
                  if ((13'sd4426/*4426:xpc10*/==xpc10))  xpc10 <= 13'sd4427/*4427:xpc10*/;
                  if ((13'sd4427/*4427:xpc10*/==xpc10))  xpc10 <= 13'sd4428/*4428:xpc10*/;
                  if ((13'sd4431/*4431:xpc10*/==xpc10))  xpc10 <= 13'sd4432/*4432:xpc10*/;
                  if ((13'sd4432/*4432:xpc10*/==xpc10))  xpc10 <= 13'sd4433/*4433:xpc10*/;
                  if ((13'sd4433/*4433:xpc10*/==xpc10))  xpc10 <= 13'sd4434/*4434:xpc10*/;
                  if ((13'sd4435/*4435:xpc10*/==xpc10))  xpc10 <= 13'sd4436/*4436:xpc10*/;
                  if ((13'sd4436/*4436:xpc10*/==xpc10))  xpc10 <= 13'sd4437/*4437:xpc10*/;
                  if ((13'sd4437/*4437:xpc10*/==xpc10))  xpc10 <= 13'sd4438/*4438:xpc10*/;
                  if ((13'sd4441/*4441:xpc10*/==xpc10))  xpc10 <= 13'sd4442/*4442:xpc10*/;
                  if ((13'sd4442/*4442:xpc10*/==xpc10))  xpc10 <= 13'sd4443/*4443:xpc10*/;
                  if ((13'sd4443/*4443:xpc10*/==xpc10))  xpc10 <= 13'sd4444/*4444:xpc10*/;
                  if ((13'sd4445/*4445:xpc10*/==xpc10))  xpc10 <= 13'sd4446/*4446:xpc10*/;
                  if ((13'sd4446/*4446:xpc10*/==xpc10))  xpc10 <= 13'sd4447/*4447:xpc10*/;
                  if ((13'sd4447/*4447:xpc10*/==xpc10))  xpc10 <= 13'sd4448/*4448:xpc10*/;
                  if ((13'sd4452/*4452:xpc10*/==xpc10))  xpc10 <= 13'sd4453/*4453:xpc10*/;
                  if ((13'sd4453/*4453:xpc10*/==xpc10))  xpc10 <= 13'sd4454/*4454:xpc10*/;
                  if ((13'sd4454/*4454:xpc10*/==xpc10))  xpc10 <= 13'sd4455/*4455:xpc10*/;
                  if ((13'sd4455/*4455:xpc10*/==xpc10))  xpc10 <= 13'sd4456/*4456:xpc10*/;
                  if ((13'sd4456/*4456:xpc10*/==xpc10))  xpc10 <= 13'sd4457/*4457:xpc10*/;
                  if ((13'sd4457/*4457:xpc10*/==xpc10))  xpc10 <= 13'sd4458/*4458:xpc10*/;
                  if ((13'sd4458/*4458:xpc10*/==xpc10))  xpc10 <= 13'sd4459/*4459:xpc10*/;
                  if ((13'sd4460/*4460:xpc10*/==xpc10))  xpc10 <= 13'sd4461/*4461:xpc10*/;
                  if ((13'sd4461/*4461:xpc10*/==xpc10))  xpc10 <= 13'sd4462/*4462:xpc10*/;
                  if ((13'sd4462/*4462:xpc10*/==xpc10))  xpc10 <= 13'sd4463/*4463:xpc10*/;
                  if ((13'sd4464/*4464:xpc10*/==xpc10))  xpc10 <= 13'sd4465/*4465:xpc10*/;
                  if ((13'sd4465/*4465:xpc10*/==xpc10))  xpc10 <= 13'sd4466/*4466:xpc10*/;
                  if ((13'sd4466/*4466:xpc10*/==xpc10))  xpc10 <= 13'sd4467/*4467:xpc10*/;
                  if ((13'sd4468/*4468:xpc10*/==xpc10))  xpc10 <= 13'sd511/*511:xpc10*/;
                  if ((13'sd4469/*4469:xpc10*/==xpc10))  xpc10 <= 13'sd4470/*4470:xpc10*/;
                  if ((13'sd4470/*4470:xpc10*/==xpc10))  xpc10 <= 13'sd4471/*4471:xpc10*/;
                  if ((13'sd4472/*4472:xpc10*/==xpc10))  xpc10 <= 13'sd4473/*4473:xpc10*/;
                  if ((13'sd4473/*4473:xpc10*/==xpc10))  xpc10 <= 13'sd4474/*4474:xpc10*/;
                  if ((13'sd4474/*4474:xpc10*/==xpc10))  xpc10 <= 13'sd4475/*4475:xpc10*/;
                  if ((13'sd4476/*4476:xpc10*/==xpc10))  xpc10 <= 13'sd4465/*4465:xpc10*/;
                  if ((13'sd4477/*4477:xpc10*/==xpc10))  xpc10 <= 13'sd4478/*4478:xpc10*/;
                  if ((13'sd4478/*4478:xpc10*/==xpc10))  xpc10 <= 13'sd4479/*4479:xpc10*/;
                  if ((13'sd4480/*4480:xpc10*/==xpc10))  xpc10 <= 13'sd4481/*4481:xpc10*/;
                  if ((13'sd4481/*4481:xpc10*/==xpc10))  xpc10 <= 13'sd4482/*4482:xpc10*/;
                  if ((13'sd4482/*4482:xpc10*/==xpc10))  xpc10 <= 13'sd4483/*4483:xpc10*/;
                  if ((13'sd4484/*4484:xpc10*/==xpc10))  xpc10 <= 13'sd4465/*4465:xpc10*/;
                  if ((13'sd4485/*4485:xpc10*/==xpc10))  xpc10 <= 13'sd4486/*4486:xpc10*/;
                  if ((13'sd4486/*4486:xpc10*/==xpc10))  xpc10 <= 13'sd4487/*4487:xpc10*/;
                  if ((13'sd4488/*4488:xpc10*/==xpc10))  xpc10 <= 13'sd4465/*4465:xpc10*/;
                  if ((13'sd4489/*4489:xpc10*/==xpc10))  xpc10 <= 13'sd4490/*4490:xpc10*/;
                  if ((13'sd4490/*4490:xpc10*/==xpc10))  xpc10 <= 13'sd4491/*4491:xpc10*/;
                  if ((13'sd4492/*4492:xpc10*/==xpc10))  xpc10 <= 13'sd4446/*4446:xpc10*/;
                  if ((13'sd4493/*4493:xpc10*/==xpc10))  xpc10 <= 13'sd4494/*4494:xpc10*/;
                  if ((13'sd4494/*4494:xpc10*/==xpc10))  xpc10 <= 13'sd4495/*4495:xpc10*/;
                  if ((13'sd4496/*4496:xpc10*/==xpc10))  xpc10 <= 13'sd4436/*4436:xpc10*/;
                  if ((13'sd4497/*4497:xpc10*/==xpc10))  xpc10 <= 13'sd4498/*4498:xpc10*/;
                  if ((13'sd4498/*4498:xpc10*/==xpc10))  xpc10 <= 13'sd4499/*4499:xpc10*/;
                  if ((13'sd4500/*4500:xpc10*/==xpc10))  xpc10 <= 13'sd4501/*4501:xpc10*/;
                  if ((13'sd4501/*4501:xpc10*/==xpc10))  xpc10 <= 13'sd4502/*4502:xpc10*/;
                  if ((13'sd4502/*4502:xpc10*/==xpc10))  xpc10 <= 13'sd4503/*4503:xpc10*/;
                  if ((13'sd4504/*4504:xpc10*/==xpc10))  xpc10 <= 13'sd4505/*4505:xpc10*/;
                  if ((13'sd4505/*4505:xpc10*/==xpc10))  xpc10 <= 13'sd4506/*4506:xpc10*/;
                  if ((13'sd4506/*4506:xpc10*/==xpc10))  xpc10 <= 13'sd4507/*4507:xpc10*/;
                  if ((13'sd4507/*4507:xpc10*/==xpc10))  xpc10 <= 13'sd4508/*4508:xpc10*/;
                  if ((13'sd4509/*4509:xpc10*/==xpc10))  xpc10 <= 13'sd511/*511:xpc10*/;
                  if ((13'sd4510/*4510:xpc10*/==xpc10))  xpc10 <= 13'sd4511/*4511:xpc10*/;
                  if ((13'sd4511/*4511:xpc10*/==xpc10))  xpc10 <= 13'sd4512/*4512:xpc10*/;
                  if ((13'sd4513/*4513:xpc10*/==xpc10))  xpc10 <= 13'sd4514/*4514:xpc10*/;
                  if ((13'sd4514/*4514:xpc10*/==xpc10))  xpc10 <= 13'sd4515/*4515:xpc10*/;
                  if ((13'sd4515/*4515:xpc10*/==xpc10))  xpc10 <= 13'sd4516/*4516:xpc10*/;
                  if ((13'sd4517/*4517:xpc10*/==xpc10))  xpc10 <= 13'sd4518/*4518:xpc10*/;
                  if ((13'sd4518/*4518:xpc10*/==xpc10))  xpc10 <= 13'sd4519/*4519:xpc10*/;
                  if ((13'sd4519/*4519:xpc10*/==xpc10))  xpc10 <= 13'sd4520/*4520:xpc10*/;
                  if ((13'sd4521/*4521:xpc10*/==xpc10))  xpc10 <= 13'sd511/*511:xpc10*/;
                  if ((13'sd4522/*4522:xpc10*/==xpc10))  xpc10 <= 13'sd4523/*4523:xpc10*/;
                  if ((13'sd4523/*4523:xpc10*/==xpc10))  xpc10 <= 13'sd4524/*4524:xpc10*/;
                  if ((13'sd4525/*4525:xpc10*/==xpc10))  xpc10 <= 13'sd4518/*4518:xpc10*/;
                  if ((13'sd4526/*4526:xpc10*/==xpc10))  xpc10 <= 13'sd4527/*4527:xpc10*/;
                  if ((13'sd4527/*4527:xpc10*/==xpc10))  xpc10 <= 13'sd4528/*4528:xpc10*/;
                  if ((13'sd4529/*4529:xpc10*/==xpc10))  xpc10 <= 13'sd4530/*4530:xpc10*/;
                  if ((13'sd4530/*4530:xpc10*/==xpc10))  xpc10 <= 13'sd4531/*4531:xpc10*/;
                  if ((13'sd4531/*4531:xpc10*/==xpc10))  xpc10 <= 13'sd4532/*4532:xpc10*/;
                  if ((13'sd4533/*4533:xpc10*/==xpc10))  xpc10 <= 13'sd4534/*4534:xpc10*/;
                  if ((13'sd4534/*4534:xpc10*/==xpc10))  xpc10 <= 13'sd4535/*4535:xpc10*/;
                  if ((13'sd4535/*4535:xpc10*/==xpc10))  xpc10 <= 13'sd4536/*4536:xpc10*/;
                  if ((13'sd4537/*4537:xpc10*/==xpc10))  xpc10 <= 13'sd4538/*4538:xpc10*/;
                  if ((13'sd4538/*4538:xpc10*/==xpc10))  xpc10 <= 13'sd4539/*4539:xpc10*/;
                  if ((13'sd4539/*4539:xpc10*/==xpc10))  xpc10 <= 13'sd4540/*4540:xpc10*/;
                  if ((13'sd4541/*4541:xpc10*/==xpc10))  xpc10 <= 13'sd4542/*4542:xpc10*/;
                  if ((13'sd4542/*4542:xpc10*/==xpc10))  xpc10 <= 13'sd4543/*4543:xpc10*/;
                  if ((13'sd4543/*4543:xpc10*/==xpc10))  xpc10 <= 13'sd4544/*4544:xpc10*/;
                  if ((13'sd4545/*4545:xpc10*/==xpc10))  xpc10 <= 13'sd511/*511:xpc10*/;
                  if ((13'sd4546/*4546:xpc10*/==xpc10))  xpc10 <= 13'sd4547/*4547:xpc10*/;
                  if ((13'sd4547/*4547:xpc10*/==xpc10))  xpc10 <= 13'sd4548/*4548:xpc10*/;
                  if ((13'sd4549/*4549:xpc10*/==xpc10))  xpc10 <= 13'sd4542/*4542:xpc10*/;
                  if ((13'sd4550/*4550:xpc10*/==xpc10))  xpc10 <= 13'sd4551/*4551:xpc10*/;
                  if ((13'sd4551/*4551:xpc10*/==xpc10))  xpc10 <= 13'sd4552/*4552:xpc10*/;
                  if ((13'sd4555/*4555:xpc10*/==xpc10))  xpc10 <= 13'sd4556/*4556:xpc10*/;
                  if ((13'sd4556/*4556:xpc10*/==xpc10))  xpc10 <= 13'sd4557/*4557:xpc10*/;
                  if ((13'sd4557/*4557:xpc10*/==xpc10))  xpc10 <= 13'sd4558/*4558:xpc10*/;
                  if ((13'sd4559/*4559:xpc10*/==xpc10))  xpc10 <= 13'sd4560/*4560:xpc10*/;
                  if ((13'sd4560/*4560:xpc10*/==xpc10))  xpc10 <= 13'sd4561/*4561:xpc10*/;
                  if ((13'sd4561/*4561:xpc10*/==xpc10))  xpc10 <= 13'sd4562/*4562:xpc10*/;
                  if ((13'sd4565/*4565:xpc10*/==xpc10))  xpc10 <= 13'sd4566/*4566:xpc10*/;
                  if ((13'sd4566/*4566:xpc10*/==xpc10))  xpc10 <= 13'sd4567/*4567:xpc10*/;
                  if ((13'sd4567/*4567:xpc10*/==xpc10))  xpc10 <= 13'sd4568/*4568:xpc10*/;
                  if ((13'sd4570/*4570:xpc10*/==xpc10))  xpc10 <= 13'sd4571/*4571:xpc10*/;
                  if ((13'sd4571/*4571:xpc10*/==xpc10))  xpc10 <= 13'sd4572/*4572:xpc10*/;
                  if ((13'sd4572/*4572:xpc10*/==xpc10))  xpc10 <= 13'sd4573/*4573:xpc10*/;
                  if ((13'sd4574/*4574:xpc10*/==xpc10))  xpc10 <= 13'sd4575/*4575:xpc10*/;
                  if ((13'sd4575/*4575:xpc10*/==xpc10))  xpc10 <= 13'sd4576/*4576:xpc10*/;
                  if ((13'sd4576/*4576:xpc10*/==xpc10))  xpc10 <= 13'sd4577/*4577:xpc10*/;
                  if ((13'sd4579/*4579:xpc10*/==xpc10))  xpc10 <= 13'sd4580/*4580:xpc10*/;
                  if ((13'sd4580/*4580:xpc10*/==xpc10))  xpc10 <= 13'sd4581/*4581:xpc10*/;
                  if ((13'sd4581/*4581:xpc10*/==xpc10))  xpc10 <= 13'sd4582/*4582:xpc10*/;
                  if ((13'sd4587/*4587:xpc10*/==xpc10))  xpc10 <= 13'sd4588/*4588:xpc10*/;
                  if ((13'sd4588/*4588:xpc10*/==xpc10))  xpc10 <= 13'sd4589/*4589:xpc10*/;
                  if ((13'sd4589/*4589:xpc10*/==xpc10))  xpc10 <= 13'sd4590/*4590:xpc10*/;
                  if ((13'sd4591/*4591:xpc10*/==xpc10))  xpc10 <= 13'sd4592/*4592:xpc10*/;
                  if ((13'sd4592/*4592:xpc10*/==xpc10))  xpc10 <= 13'sd4593/*4593:xpc10*/;
                  if ((13'sd4593/*4593:xpc10*/==xpc10))  xpc10 <= 13'sd4594/*4594:xpc10*/;
                  if ((13'sd4595/*4595:xpc10*/==xpc10))  xpc10 <= 13'sd4596/*4596:xpc10*/;
                  if ((13'sd4596/*4596:xpc10*/==xpc10))  xpc10 <= 13'sd4597/*4597:xpc10*/;
                  if ((13'sd4597/*4597:xpc10*/==xpc10))  xpc10 <= 13'sd4598/*4598:xpc10*/;
                  if ((13'sd4599/*4599:xpc10*/==xpc10))  xpc10 <= 13'sd4600/*4600:xpc10*/;
                  if ((13'sd4600/*4600:xpc10*/==xpc10))  xpc10 <= 13'sd4601/*4601:xpc10*/;
                  if ((13'sd4601/*4601:xpc10*/==xpc10))  xpc10 <= 13'sd4602/*4602:xpc10*/;
                  if ((13'sd4603/*4603:xpc10*/==xpc10))  xpc10 <= 13'sd4604/*4604:xpc10*/;
                  if ((13'sd4604/*4604:xpc10*/==xpc10))  xpc10 <= 13'sd4605/*4605:xpc10*/;
                  if ((13'sd4605/*4605:xpc10*/==xpc10))  xpc10 <= 13'sd4606/*4606:xpc10*/;
                  if ((13'sd4607/*4607:xpc10*/==xpc10))  xpc10 <= 13'sd511/*511:xpc10*/;
                  if ((13'sd4608/*4608:xpc10*/==xpc10))  xpc10 <= 13'sd4609/*4609:xpc10*/;
                  if ((13'sd4609/*4609:xpc10*/==xpc10))  xpc10 <= 13'sd4610/*4610:xpc10*/;
                  if ((13'sd4611/*4611:xpc10*/==xpc10))  xpc10 <= 13'sd4604/*4604:xpc10*/;
                  if ((13'sd4612/*4612:xpc10*/==xpc10))  xpc10 <= 13'sd4613/*4613:xpc10*/;
                  if ((13'sd4613/*4613:xpc10*/==xpc10))  xpc10 <= 13'sd4614/*4614:xpc10*/;
                  if ((13'sd4617/*4617:xpc10*/==xpc10))  xpc10 <= 13'sd4618/*4618:xpc10*/;
                  if ((13'sd4618/*4618:xpc10*/==xpc10))  xpc10 <= 13'sd4619/*4619:xpc10*/;
                  if ((13'sd4619/*4619:xpc10*/==xpc10))  xpc10 <= 13'sd4620/*4620:xpc10*/;
                  if ((13'sd4621/*4621:xpc10*/==xpc10))  xpc10 <= 13'sd4622/*4622:xpc10*/;
                  if ((13'sd4622/*4622:xpc10*/==xpc10))  xpc10 <= 13'sd4623/*4623:xpc10*/;
                  if ((13'sd4623/*4623:xpc10*/==xpc10))  xpc10 <= 13'sd4624/*4624:xpc10*/;
                  if ((13'sd4627/*4627:xpc10*/==xpc10))  xpc10 <= 13'sd4628/*4628:xpc10*/;
                  if ((13'sd4628/*4628:xpc10*/==xpc10))  xpc10 <= 13'sd4629/*4629:xpc10*/;
                  if ((13'sd4629/*4629:xpc10*/==xpc10))  xpc10 <= 13'sd4630/*4630:xpc10*/;
                  if ((13'sd4632/*4632:xpc10*/==xpc10))  xpc10 <= 13'sd4633/*4633:xpc10*/;
                  if ((13'sd4633/*4633:xpc10*/==xpc10))  xpc10 <= 13'sd4634/*4634:xpc10*/;
                  if ((13'sd4634/*4634:xpc10*/==xpc10))  xpc10 <= 13'sd4635/*4635:xpc10*/;
                  if ((13'sd4636/*4636:xpc10*/==xpc10))  xpc10 <= 13'sd4637/*4637:xpc10*/;
                  if ((13'sd4637/*4637:xpc10*/==xpc10))  xpc10 <= 13'sd4638/*4638:xpc10*/;
                  if ((13'sd4638/*4638:xpc10*/==xpc10))  xpc10 <= 13'sd4639/*4639:xpc10*/;
                  if ((13'sd4641/*4641:xpc10*/==xpc10))  xpc10 <= 13'sd4642/*4642:xpc10*/;
                  if ((13'sd4642/*4642:xpc10*/==xpc10))  xpc10 <= 13'sd4643/*4643:xpc10*/;
                  if ((13'sd4643/*4643:xpc10*/==xpc10))  xpc10 <= 13'sd4644/*4644:xpc10*/;
                  if ((13'sd4649/*4649:xpc10*/==xpc10))  xpc10 <= 13'sd4650/*4650:xpc10*/;
                  if ((13'sd4650/*4650:xpc10*/==xpc10))  xpc10 <= 13'sd4651/*4651:xpc10*/;
                  if ((13'sd4651/*4651:xpc10*/==xpc10))  xpc10 <= 13'sd4652/*4652:xpc10*/;
                  if ((13'sd4665/*4665:xpc10*/==xpc10))  xpc10 <= 13'sd4666/*4666:xpc10*/;
                  if ((13'sd4666/*4666:xpc10*/==xpc10))  xpc10 <= 13'sd4667/*4667:xpc10*/;
                  if ((13'sd4667/*4667:xpc10*/==xpc10))  xpc10 <= 13'sd4668/*4668:xpc10*/;
                  if ((13'sd4668/*4668:xpc10*/==xpc10))  xpc10 <= 13'sd4669/*4669:xpc10*/;
                  if ((13'sd4669/*4669:xpc10*/==xpc10))  xpc10 <= 13'sd4670/*4670:xpc10*/;
                  if ((13'sd4670/*4670:xpc10*/==xpc10))  xpc10 <= 13'sd4671/*4671:xpc10*/;
                  if ((13'sd4671/*4671:xpc10*/==xpc10))  xpc10 <= 13'sd4672/*4672:xpc10*/;
                  if ((13'sd4672/*4672:xpc10*/==xpc10))  xpc10 <= 13'sd4673/*4673:xpc10*/;
                  if ((13'sd4677/*4677:xpc10*/==xpc10))  xpc10 <= 13'sd4678/*4678:xpc10*/;
                  if ((13'sd4678/*4678:xpc10*/==xpc10))  xpc10 <= 13'sd4679/*4679:xpc10*/;
                  if ((13'sd4679/*4679:xpc10*/==xpc10))  xpc10 <= 13'sd4680/*4680:xpc10*/;
                  if ((13'sd4682/*4682:xpc10*/==xpc10))  xpc10 <= 13'sd4683/*4683:xpc10*/;
                  if ((13'sd4683/*4683:xpc10*/==xpc10))  xpc10 <= 13'sd4684/*4684:xpc10*/;
                  if ((13'sd4684/*4684:xpc10*/==xpc10))  xpc10 <= 13'sd4685/*4685:xpc10*/;
                  if ((13'sd4692/*4692:xpc10*/==xpc10))  xpc10 <= 13'sd4693/*4693:xpc10*/;
                  if ((13'sd4693/*4693:xpc10*/==xpc10))  xpc10 <= 13'sd4694/*4694:xpc10*/;
                  if ((13'sd4694/*4694:xpc10*/==xpc10))  xpc10 <= 13'sd4695/*4695:xpc10*/;
                  if ((13'sd4697/*4697:xpc10*/==xpc10))  xpc10 <= 13'sd4698/*4698:xpc10*/;
                  if ((13'sd4698/*4698:xpc10*/==xpc10))  xpc10 <= 13'sd4699/*4699:xpc10*/;
                  if ((13'sd4699/*4699:xpc10*/==xpc10))  xpc10 <= 13'sd4700/*4700:xpc10*/;
                  if ((13'sd4707/*4707:xpc10*/==xpc10))  xpc10 <= 13'sd4708/*4708:xpc10*/;
                  if ((13'sd4708/*4708:xpc10*/==xpc10))  xpc10 <= 13'sd4709/*4709:xpc10*/;
                  if ((13'sd4709/*4709:xpc10*/==xpc10))  xpc10 <= 13'sd4710/*4710:xpc10*/;
                  if ((13'sd4712/*4712:xpc10*/==xpc10))  xpc10 <= 13'sd4713/*4713:xpc10*/;
                  if ((13'sd4713/*4713:xpc10*/==xpc10))  xpc10 <= 13'sd4714/*4714:xpc10*/;
                  if ((13'sd4714/*4714:xpc10*/==xpc10))  xpc10 <= 13'sd4715/*4715:xpc10*/;
                  if ((13'sd4717/*4717:xpc10*/==xpc10))  xpc10 <= 13'sd4718/*4718:xpc10*/;
                  if ((13'sd4718/*4718:xpc10*/==xpc10))  xpc10 <= 13'sd4719/*4719:xpc10*/;
                  if ((13'sd4719/*4719:xpc10*/==xpc10))  xpc10 <= 13'sd4720/*4720:xpc10*/;
                  if ((13'sd4722/*4722:xpc10*/==xpc10))  xpc10 <= 13'sd4723/*4723:xpc10*/;
                  if ((13'sd4723/*4723:xpc10*/==xpc10))  xpc10 <= 13'sd4724/*4724:xpc10*/;
                  if ((13'sd4724/*4724:xpc10*/==xpc10))  xpc10 <= 13'sd4725/*4725:xpc10*/;
                  if ((13'sd4727/*4727:xpc10*/==xpc10))  xpc10 <= 13'sd4728/*4728:xpc10*/;
                  if ((13'sd4728/*4728:xpc10*/==xpc10))  xpc10 <= 13'sd4729/*4729:xpc10*/;
                  if ((13'sd4730/*4730:xpc10*/==xpc10))  xpc10 <= 13'sd4731/*4731:xpc10*/;
                  if ((13'sd4731/*4731:xpc10*/==xpc10))  xpc10 <= 13'sd4732/*4732:xpc10*/;
                  if ((13'sd4732/*4732:xpc10*/==xpc10))  xpc10 <= 13'sd4733/*4733:xpc10*/;
                  if ((13'sd4735/*4735:xpc10*/==xpc10))  xpc10 <= 13'sd4736/*4736:xpc10*/;
                  if ((13'sd4736/*4736:xpc10*/==xpc10))  xpc10 <= 13'sd4737/*4737:xpc10*/;
                  if ((13'sd4737/*4737:xpc10*/==xpc10))  xpc10 <= 13'sd4738/*4738:xpc10*/;
                  if ((13'sd4739/*4739:xpc10*/==xpc10))  xpc10 <= 13'sd4740/*4740:xpc10*/;
                  if ((13'sd4740/*4740:xpc10*/==xpc10))  xpc10 <= 13'sd4741/*4741:xpc10*/;
                  if ((13'sd4741/*4741:xpc10*/==xpc10))  xpc10 <= 13'sd4742/*4742:xpc10*/;
                  if ((13'sd4743/*4743:xpc10*/==xpc10))  xpc10 <= 13'sd4744/*4744:xpc10*/;
                  if ((13'sd4744/*4744:xpc10*/==xpc10))  xpc10 <= 13'sd4745/*4745:xpc10*/;
                  if ((13'sd4745/*4745:xpc10*/==xpc10))  xpc10 <= 13'sd4746/*4746:xpc10*/;
                  if ((13'sd4747/*4747:xpc10*/==xpc10))  xpc10 <= 13'sd4748/*4748:xpc10*/;
                  if ((13'sd4748/*4748:xpc10*/==xpc10))  xpc10 <= 13'sd4749/*4749:xpc10*/;
                  if ((13'sd4749/*4749:xpc10*/==xpc10))  xpc10 <= 13'sd4750/*4750:xpc10*/;
                  if ((13'sd4750/*4750:xpc10*/==xpc10))  xpc10 <= 13'sd4751/*4751:xpc10*/;
                  if ((13'sd4752/*4752:xpc10*/==xpc10))  xpc10 <= 13'sd4753/*4753:xpc10*/;
                  if ((13'sd4753/*4753:xpc10*/==xpc10))  xpc10 <= 13'sd4754/*4754:xpc10*/;
                  if ((13'sd4754/*4754:xpc10*/==xpc10))  xpc10 <= 13'sd4755/*4755:xpc10*/;
                  if ((13'sd4756/*4756:xpc10*/==xpc10))  xpc10 <= 13'sd4757/*4757:xpc10*/;
                  if ((13'sd4757/*4757:xpc10*/==xpc10))  xpc10 <= 13'sd4758/*4758:xpc10*/;
                  if ((13'sd4758/*4758:xpc10*/==xpc10))  xpc10 <= 13'sd4759/*4759:xpc10*/;
                  if ((13'sd4763/*4763:xpc10*/==xpc10))  xpc10 <= 13'sd4764/*4764:xpc10*/;
                  if ((13'sd4764/*4764:xpc10*/==xpc10))  xpc10 <= 13'sd4765/*4765:xpc10*/;
                  if ((13'sd4765/*4765:xpc10*/==xpc10))  xpc10 <= 13'sd4766/*4766:xpc10*/;
                  if ((13'sd4768/*4768:xpc10*/==xpc10))  xpc10 <= 13'sd4769/*4769:xpc10*/;
                  if ((13'sd4769/*4769:xpc10*/==xpc10))  xpc10 <= 13'sd4770/*4770:xpc10*/;
                  if ((13'sd4770/*4770:xpc10*/==xpc10))  xpc10 <= 13'sd4771/*4771:xpc10*/;
                  if ((13'sd4772/*4772:xpc10*/==xpc10))  xpc10 <= 13'sd4773/*4773:xpc10*/;
                  if ((13'sd4773/*4773:xpc10*/==xpc10))  xpc10 <= 13'sd4774/*4774:xpc10*/;
                  if ((13'sd4774/*4774:xpc10*/==xpc10))  xpc10 <= 13'sd4775/*4775:xpc10*/;
                  if ((13'sd4776/*4776:xpc10*/==xpc10))  xpc10 <= 13'sd511/*511:xpc10*/;
                  if ((13'sd4777/*4777:xpc10*/==xpc10))  xpc10 <= 13'sd4778/*4778:xpc10*/;
                  if ((13'sd4778/*4778:xpc10*/==xpc10))  xpc10 <= 13'sd4779/*4779:xpc10*/;
                  if ((13'sd4781/*4781:xpc10*/==xpc10))  xpc10 <= 13'sd4769/*4769:xpc10*/;
                  if ((13'sd4782/*4782:xpc10*/==xpc10))  xpc10 <= 13'sd4783/*4783:xpc10*/;
                  if ((13'sd4783/*4783:xpc10*/==xpc10))  xpc10 <= 13'sd4784/*4784:xpc10*/;
                  if ((13'sd4785/*4785:xpc10*/==xpc10))  xpc10 <= 13'sd4757/*4757:xpc10*/;
                  if ((13'sd4786/*4786:xpc10*/==xpc10))  xpc10 <= 13'sd4787/*4787:xpc10*/;
                  if ((13'sd4787/*4787:xpc10*/==xpc10))  xpc10 <= 13'sd4788/*4788:xpc10*/;
                  if ((13'sd4789/*4789:xpc10*/==xpc10))  xpc10 <= 13'sd4790/*4790:xpc10*/;
                  if ((13'sd4790/*4790:xpc10*/==xpc10))  xpc10 <= 13'sd4791/*4791:xpc10*/;
                  if ((13'sd4791/*4791:xpc10*/==xpc10))  xpc10 <= 13'sd4792/*4792:xpc10*/;
                  if ((13'sd4792/*4792:xpc10*/==xpc10))  xpc10 <= 13'sd4793/*4793:xpc10*/;
                  if ((13'sd4794/*4794:xpc10*/==xpc10))  xpc10 <= 13'sd4795/*4795:xpc10*/;
                  if ((13'sd4795/*4795:xpc10*/==xpc10))  xpc10 <= 13'sd4796/*4796:xpc10*/;
                  if ((13'sd4796/*4796:xpc10*/==xpc10))  xpc10 <= 13'sd4797/*4797:xpc10*/;
                  if ((13'sd4798/*4798:xpc10*/==xpc10))  xpc10 <= 13'sd4799/*4799:xpc10*/;
                  if ((13'sd4799/*4799:xpc10*/==xpc10))  xpc10 <= 13'sd4800/*4800:xpc10*/;
                  if ((13'sd4800/*4800:xpc10*/==xpc10))  xpc10 <= 13'sd4801/*4801:xpc10*/;
                  if ((13'sd4804/*4804:xpc10*/==xpc10))  xpc10 <= 13'sd4805/*4805:xpc10*/;
                  if ((13'sd4805/*4805:xpc10*/==xpc10))  xpc10 <= 13'sd4806/*4806:xpc10*/;
                  if ((13'sd4806/*4806:xpc10*/==xpc10))  xpc10 <= 13'sd4807/*4807:xpc10*/;
                  if ((13'sd4808/*4808:xpc10*/==xpc10))  xpc10 <= 13'sd4809/*4809:xpc10*/;
                  if ((13'sd4809/*4809:xpc10*/==xpc10))  xpc10 <= 13'sd4810/*4810:xpc10*/;
                  if ((13'sd4810/*4810:xpc10*/==xpc10))  xpc10 <= 13'sd4811/*4811:xpc10*/;
                  if ((13'sd4811/*4811:xpc10*/==xpc10))  xpc10 <= 13'sd4812/*4812:xpc10*/;
                  if ((13'sd4812/*4812:xpc10*/==xpc10))  xpc10 <= 13'sd4813/*4813:xpc10*/;
                  if ((13'sd4813/*4813:xpc10*/==xpc10))  xpc10 <= 13'sd4814/*4814:xpc10*/;
                  if ((13'sd4814/*4814:xpc10*/==xpc10))  xpc10 <= 13'sd4815/*4815:xpc10*/;
                  if ((13'sd4816/*4816:xpc10*/==xpc10))  xpc10 <= 13'sd4817/*4817:xpc10*/;
                  if ((13'sd4817/*4817:xpc10*/==xpc10))  xpc10 <= 13'sd4818/*4818:xpc10*/;
                  if ((13'sd4818/*4818:xpc10*/==xpc10))  xpc10 <= 13'sd4819/*4819:xpc10*/;
                  if ((13'sd4819/*4819:xpc10*/==xpc10))  xpc10 <= 13'sd4820/*4820:xpc10*/;
                  if ((13'sd4820/*4820:xpc10*/==xpc10))  xpc10 <= 13'sd4821/*4821:xpc10*/;
                  if ((13'sd4821/*4821:xpc10*/==xpc10))  xpc10 <= 13'sd4822/*4822:xpc10*/;
                  if ((13'sd4822/*4822:xpc10*/==xpc10))  xpc10 <= 13'sd4823/*4823:xpc10*/;
                  if ((13'sd4825/*4825:xpc10*/==xpc10))  xpc10 <= 13'sd4826/*4826:xpc10*/;
                  if ((13'sd4826/*4826:xpc10*/==xpc10))  xpc10 <= 13'sd4827/*4827:xpc10*/;
                  if ((13'sd4827/*4827:xpc10*/==xpc10))  xpc10 <= 13'sd4828/*4828:xpc10*/;
                  if ((13'sd4829/*4829:xpc10*/==xpc10))  xpc10 <= 13'sd4830/*4830:xpc10*/;
                  if ((13'sd4830/*4830:xpc10*/==xpc10))  xpc10 <= 13'sd4831/*4831:xpc10*/;
                  if ((13'sd4831/*4831:xpc10*/==xpc10))  xpc10 <= 13'sd4832/*4832:xpc10*/;
                  if ((13'sd4833/*4833:xpc10*/==xpc10))  xpc10 <= 13'sd4834/*4834:xpc10*/;
                  if ((13'sd4834/*4834:xpc10*/==xpc10))  xpc10 <= 13'sd4835/*4835:xpc10*/;
                  if ((13'sd4835/*4835:xpc10*/==xpc10))  xpc10 <= 13'sd4836/*4836:xpc10*/;
                  if ((13'sd4837/*4837:xpc10*/==xpc10))  xpc10 <= 13'sd4838/*4838:xpc10*/;
                  if ((13'sd4838/*4838:xpc10*/==xpc10))  xpc10 <= 13'sd4839/*4839:xpc10*/;
                  if ((13'sd4839/*4839:xpc10*/==xpc10))  xpc10 <= 13'sd4840/*4840:xpc10*/;
                  if ((13'sd4841/*4841:xpc10*/==xpc10))  xpc10 <= 13'sd4842/*4842:xpc10*/;
                  if ((13'sd4842/*4842:xpc10*/==xpc10))  xpc10 <= 13'sd4843/*4843:xpc10*/;
                  if ((13'sd4843/*4843:xpc10*/==xpc10))  xpc10 <= 13'sd4844/*4844:xpc10*/;
                  if ((13'sd4845/*4845:xpc10*/==xpc10))  xpc10 <= 13'sd4846/*4846:xpc10*/;
                  if ((13'sd4846/*4846:xpc10*/==xpc10))  xpc10 <= 13'sd4847/*4847:xpc10*/;
                  if ((13'sd4847/*4847:xpc10*/==xpc10))  xpc10 <= 13'sd4848/*4848:xpc10*/;
                  if ((13'sd4849/*4849:xpc10*/==xpc10))  xpc10 <= 13'sd4773/*4773:xpc10*/;
                  if ((13'sd4850/*4850:xpc10*/==xpc10))  xpc10 <= 13'sd4851/*4851:xpc10*/;
                  if ((13'sd4851/*4851:xpc10*/==xpc10))  xpc10 <= 13'sd4852/*4852:xpc10*/;
                  if ((13'sd4853/*4853:xpc10*/==xpc10))  xpc10 <= 13'sd4846/*4846:xpc10*/;
                  if ((13'sd4854/*4854:xpc10*/==xpc10))  xpc10 <= 13'sd4855/*4855:xpc10*/;
                  if ((13'sd4855/*4855:xpc10*/==xpc10))  xpc10 <= 13'sd4856/*4856:xpc10*/;
                  if ((13'sd4857/*4857:xpc10*/==xpc10))  xpc10 <= 13'sd4858/*4858:xpc10*/;
                  if ((13'sd4858/*4858:xpc10*/==xpc10))  xpc10 <= 13'sd4859/*4859:xpc10*/;
                  if ((13'sd4859/*4859:xpc10*/==xpc10))  xpc10 <= 13'sd4860/*4860:xpc10*/;
                  if ((13'sd4864/*4864:xpc10*/==xpc10))  xpc10 <= 13'sd4865/*4865:xpc10*/;
                  if ((13'sd4865/*4865:xpc10*/==xpc10))  xpc10 <= 13'sd4866/*4866:xpc10*/;
                  if ((13'sd4866/*4866:xpc10*/==xpc10))  xpc10 <= 13'sd4867/*4867:xpc10*/;
                  if ((13'sd4869/*4869:xpc10*/==xpc10))  xpc10 <= 13'sd4870/*4870:xpc10*/;
                  if ((13'sd4870/*4870:xpc10*/==xpc10))  xpc10 <= 13'sd4871/*4871:xpc10*/;
                  if ((13'sd4871/*4871:xpc10*/==xpc10))  xpc10 <= 13'sd4872/*4872:xpc10*/;
                  if ((13'sd4873/*4873:xpc10*/==xpc10))  xpc10 <= 13'sd4799/*4799:xpc10*/;
                  if ((13'sd4874/*4874:xpc10*/==xpc10))  xpc10 <= 13'sd4875/*4875:xpc10*/;
                  if ((13'sd4875/*4875:xpc10*/==xpc10))  xpc10 <= 13'sd4876/*4876:xpc10*/;
                  if ((13'sd4878/*4878:xpc10*/==xpc10))  xpc10 <= 13'sd4870/*4870:xpc10*/;
                  if ((13'sd4879/*4879:xpc10*/==xpc10))  xpc10 <= 13'sd4880/*4880:xpc10*/;
                  if ((13'sd4880/*4880:xpc10*/==xpc10))  xpc10 <= 13'sd4881/*4881:xpc10*/;
                  if ((13'sd4882/*4882:xpc10*/==xpc10))  xpc10 <= 13'sd4883/*4883:xpc10*/;
                  if ((13'sd4883/*4883:xpc10*/==xpc10))  xpc10 <= 13'sd4884/*4884:xpc10*/;
                  if ((13'sd4884/*4884:xpc10*/==xpc10))  xpc10 <= 13'sd4885/*4885:xpc10*/;
                  if ((13'sd4886/*4886:xpc10*/==xpc10))  xpc10 <= 13'sd4887/*4887:xpc10*/;
                  if ((13'sd4887/*4887:xpc10*/==xpc10))  xpc10 <= 13'sd4888/*4888:xpc10*/;
                  if ((13'sd4888/*4888:xpc10*/==xpc10))  xpc10 <= 13'sd4889/*4889:xpc10*/;
                  if ((13'sd4890/*4890:xpc10*/==xpc10))  xpc10 <= 13'sd4799/*4799:xpc10*/;
                  if ((13'sd4891/*4891:xpc10*/==xpc10))  xpc10 <= 13'sd4892/*4892:xpc10*/;
                  if ((13'sd4892/*4892:xpc10*/==xpc10))  xpc10 <= 13'sd4893/*4893:xpc10*/;
                  if ((13'sd4894/*4894:xpc10*/==xpc10))  xpc10 <= 13'sd4887/*4887:xpc10*/;
                  if ((13'sd4895/*4895:xpc10*/==xpc10))  xpc10 <= 13'sd4896/*4896:xpc10*/;
                  if ((13'sd4896/*4896:xpc10*/==xpc10))  xpc10 <= 13'sd4897/*4897:xpc10*/;
                  if ((13'sd4899/*4899:xpc10*/==xpc10))  xpc10 <= 13'sd4713/*4713:xpc10*/;
                  if ((13'sd4900/*4900:xpc10*/==xpc10))  xpc10 <= 13'sd4901/*4901:xpc10*/;
                  if ((13'sd4901/*4901:xpc10*/==xpc10))  xpc10 <= 13'sd4902/*4902:xpc10*/;
                  if ((13'sd4904/*4904:xpc10*/==xpc10))  xpc10 <= 13'sd4698/*4698:xpc10*/;
                  if ((13'sd4905/*4905:xpc10*/==xpc10))  xpc10 <= 13'sd4906/*4906:xpc10*/;
                  if ((13'sd4906/*4906:xpc10*/==xpc10))  xpc10 <= 13'sd4907/*4907:xpc10*/;
                  if ((13'sd4909/*4909:xpc10*/==xpc10))  xpc10 <= 13'sd4683/*4683:xpc10*/;
                  if ((13'sd4910/*4910:xpc10*/==xpc10))  xpc10 <= 13'sd4911/*4911:xpc10*/;
                  if ((13'sd4911/*4911:xpc10*/==xpc10))  xpc10 <= 13'sd4912/*4912:xpc10*/;
                  if ((13'sd4912/*4912:xpc10*/==xpc10))  xpc10 <= 13'sd4913/*4913:xpc10*/;
                  if ((13'sd4913/*4913:xpc10*/==xpc10))  xpc10 <= 13'sd4670/*4670:xpc10*/;
                  if ((13'sd4914/*4914:xpc10*/==xpc10))  xpc10 <= 13'sd4915/*4915:xpc10*/;
                  if ((13'sd4915/*4915:xpc10*/==xpc10))  xpc10 <= 13'sd4916/*4916:xpc10*/;
                  if ((13'sd4917/*4917:xpc10*/==xpc10))  xpc10 <= 13'sd4622/*4622:xpc10*/;
                  if ((13'sd4918/*4918:xpc10*/==xpc10))  xpc10 <= 13'sd4919/*4919:xpc10*/;
                  if ((13'sd4919/*4919:xpc10*/==xpc10))  xpc10 <= 13'sd4920/*4920:xpc10*/;
                  if ((13'sd4921/*4921:xpc10*/==xpc10))  xpc10 <= 13'sd4560/*4560:xpc10*/;
                  if ((13'sd4922/*4922:xpc10*/==xpc10))  xpc10 <= 13'sd4923/*4923:xpc10*/;
                  if ((13'sd4923/*4923:xpc10*/==xpc10))  xpc10 <= 13'sd4924/*4924:xpc10*/;
                  if ((13'sd4925/*4925:xpc10*/==xpc10))  xpc10 <= 13'sd450/*450:xpc10*/;
                  if ((13'sd4926/*4926:xpc10*/==xpc10))  xpc10 <= 13'sd4927/*4927:xpc10*/;
                  if ((13'sd4927/*4927:xpc10*/==xpc10))  xpc10 <= 13'sd4928/*4928:xpc10*/;
                  if ((13'sd4929/*4929:xpc10*/==xpc10))  xpc10 <= 13'sd439/*439:xpc10*/;
                   end 
              //End structure HPR dfsin


       end 
      

// 1 vectors of width 13
// 261 vectors of width 64
// 52 vectors of width 1
// 30 vectors of width 16
// 16 vectors of width 32
// 3 vectors of width 8
// 72 array locations of width 64
// 259 array locations of width 8
// 1024 bits in scalar variables
// Total state bits in module = 25489 bits.
// Total number of leaf cells = 0
endmodule

//  
// LCP delay estimations included: turn off with -vnl-lcp-delay-estimate=disable
//HPR L/S (orangepath) auxiliary reports.
//KiwiC compilation report
//Kiwi Scientific Acceleration (KiwiC .net/CIL/C# to Verilog/SystemC compiler): Version alpha 0.2.16f : 22nd-September-2016
//23/09/2016 20:03:19
//Cmd line args:  /home/djg11/d320/hprls/kiwipro/kiwic/distro/lib/kiwic.exe -vnl-resets=synchronous -restructure2=disable -vnl-roundtrip=disable -kiwic-cil-dump=combined -kiwic-kcode-dump=enable -bevelab-default-pause-mode=maximal -bevelab-soft-pause-threshold=10 dfsin.exe ../softfloat.dll


//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation KiKiwi for prefix KiwiSystem/Kiwi

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation SyBitConverter for prefix System/BitConverter

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation CS0.4 for prefix CS/0.4

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation @8 for prefix @/8

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation CS0.2 for prefix CS/0.2

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation CS0.8 for prefix CS/0.8

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation CS0.14 for prefix CS/0.14

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation @64 for prefix @/64

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tdb0._SPILL for prefix T404/dfsin/bm_main/0.3/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tdbm0.3 for prefix T404/dfsin/bm_main/0.3

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tdsi1.5 for prefix T404/dfsin/sin/1.5

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsf0._SPILL for prefix T404/softfloat/float64_mul/0.9/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsfl0.9 for prefix T404/softfloat/float64_mul/0.9

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tse0._SPILL for prefix T404/softfloat/extractFloat64Sign/0.14/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tse0SPILL10 for prefix T404/softfloat/extractFloat64Sign/0.23/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsp4._SPILL for prefix T404/softfloat/propagateFloat64NaN/4.3/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tspr4.3 for prefix T404/softfloat/propagateFloat64NaN/4.3

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsf0SPILL10 for prefix T404/softfloat/float64_is_signaling_nan/0.6/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsf0SPILL12 for prefix T404/softfloat/float64_is_signaling_nan/0.12/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsp8._SPILL for prefix T404/softfloat/packFloat64/8.5/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsp11_SPILL for prefix T404/softfloat/propagateFloat64NaN/11.2/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tspr11.2 for prefix T404/softfloat/propagateFloat64NaN/11.2

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsp15_SPILL for prefix T404/softfloat/packFloat64/15.5/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsp18_SPILL for prefix T404/softfloat/packFloat64/18.4/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsno19.4 for prefix T404/softfloat/normalizeFloat64Subnormal/19.4

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsco0.2 for prefix T404/softfloat/countLeadingZeros64/0.2

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsco3.7 for prefix T404/softfloat/countLeadingZeros32/3.7

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsp22_SPILL for prefix T404/softfloat/packFloat64/22.4/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsno23.4 for prefix T404/softfloat/normalizeFloat64Subnormal/23.4

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsm24_SPILL for prefix T404/softfloat/mul64To128/24.24/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsmu24.24 for prefix T404/softfloat/mul64To128/24.24

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsr29_SPILL for prefix T404/softfloat/roundAndPackFloat64/29.4/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsro29.4 for prefix T404/softfloat/roundAndPackFloat64/29.4

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsp13_SPILL for prefix T404/softfloat/packFloat64/13.7/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tss18_SPILL for prefix T404/softfloat/shift64RightJamming/18.7/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tssh18.7 for prefix T404/softfloat/shift64RightJamming/18.7

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsp27_SPILL for prefix T404/softfloat/packFloat64/27.4/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsfl0.10 for prefix T404/softfloat/float64_neg/0.10

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsf1._SPILL for prefix T404/softfloat/float64_mul/1.8/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsfl1.8 for prefix T404/softfloat/float64_mul/1.8

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsi1._SPILL for prefix T404/softfloat/int32_to_float64/1.19/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsin1.19 for prefix T404/softfloat/int32_to_float64/1.19

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsco5.4 for prefix T404/softfloat/countLeadingZeros32/5.4

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsp5._SPILL for prefix T404/softfloat/packFloat64/5.21/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsf1SPILL10 for prefix T404/softfloat/float64_mul/1.24/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsfl1.24 for prefix T404/softfloat/float64_mul/1.24

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsi1SPILL10 for prefix T404/softfloat/int32_to_float64/1.34/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsin1.34 for prefix T404/softfloat/int32_to_float64/1.34

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsf1SPILL12 for prefix T404/softfloat/float64_div/1.35/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsfl1.35 for prefix T404/softfloat/float64_div/1.35

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tse0SPILL12 for prefix T404/softfloat/extractFloat64Sign/0.8/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tse0SPILL14 for prefix T404/softfloat/extractFloat64Sign/0.17/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsp2._SPILL for prefix T404/softfloat/propagateFloat64NaN/2.2/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tspr2.2 for prefix T404/softfloat/propagateFloat64NaN/2.2

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsp5SPILL10 for prefix T404/softfloat/propagateFloat64NaN/5.2/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tspr5.2 for prefix T404/softfloat/propagateFloat64NaN/5.2

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsp7._SPILL for prefix T404/softfloat/packFloat64/7.5/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsp10_SPILL for prefix T404/softfloat/propagateFloat64NaN/10.2/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tspr10.2 for prefix T404/softfloat/propagateFloat64NaN/10.2

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsp11SPILL10 for prefix T404/softfloat/packFloat64/11.5/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsp17_SPILL for prefix T404/softfloat/packFloat64/17.7/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsno18.4 for prefix T404/softfloat/normalizeFloat64Subnormal/18.4

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsp21_SPILL for prefix T404/softfloat/packFloat64/21.4/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsno22.4 for prefix T404/softfloat/normalizeFloat64Subnormal/22.4

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tse25_SPILL for prefix T404/softfloat/estimateDiv128To64/25.5/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tses25.5 for prefix T404/softfloat/estimateDiv128To64/25.5

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsm5._SPILL for prefix T404/softfloat/mul64To128/5.7/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsmu5.7 for prefix T404/softfloat/mul64To128/5.7

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tss5._SPILL for prefix T404/softfloat/sub128/5.14/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsa6._SPILL for prefix T404/softfloat/add128/6.15/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsad6.15 for prefix T404/softfloat/add128/6.15

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsm26_SPILL for prefix T404/softfloat/mul64To128/26.4/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsmu26.4 for prefix T404/softfloat/mul64To128/26.4

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tss26_SPILL for prefix T404/softfloat/sub128/26.12/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsa27_SPILL for prefix T404/softfloat/add128/27.13/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsad27.13 for prefix T404/softfloat/add128/27.13

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsr33_SPILL for prefix T404/softfloat/roundAndPackFloat64/33.4/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsro33.4 for prefix T404/softfloat/roundAndPackFloat64/33.4

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsf1SPILL14 for prefix T404/softfloat/float64_add/1.39/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsfl1.39 for prefix T404/softfloat/float64_add/1.39

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tse0SPILL16 for prefix T404/softfloat/extractFloat64Sign/0.2/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tse0SPILL18 for prefix T404/softfloat/extractFloat64Sign/0.5/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsa1._SPILL for prefix T404/softfloat/addFloat64Sigs/1.3/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsad1.3 for prefix T404/softfloat/addFloat64Sigs/1.3

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsp3._SPILL for prefix T404/softfloat/propagateFloat64NaN/3.2/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tspr3.2 for prefix T404/softfloat/propagateFloat64NaN/3.2

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tss8._SPILL for prefix T404/softfloat/shift64RightJamming/8.5/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tssh8.5 for prefix T404/softfloat/shift64RightJamming/8.5

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsp12_SPILL for prefix T404/softfloat/propagateFloat64NaN/12.2/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tspr12.2 for prefix T404/softfloat/propagateFloat64NaN/12.2

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsp13SPILL10 for prefix T404/softfloat/packFloat64/13.5/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tss17_SPILL for prefix T404/softfloat/shift64RightJamming/17.6/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tssh17.6 for prefix T404/softfloat/shift64RightJamming/17.6

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsp21SPILL10 for prefix T404/softfloat/propagateFloat64NaN/21.3/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tspr21.3 for prefix T404/softfloat/propagateFloat64NaN/21.3

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsp24_SPILL for prefix T404/softfloat/packFloat64/24.7/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsr28_SPILL for prefix T404/softfloat/roundAndPackFloat64/28.4/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsro28.4 for prefix T404/softfloat/roundAndPackFloat64/28.4

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tss2._SPILL for prefix T404/softfloat/subFloat64Sigs/2.4/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tssu2.4 for prefix T404/softfloat/subFloat64Sigs/2.4

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsp7SPILL10 for prefix T404/softfloat/propagateFloat64NaN/7.3/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tspr7.3 for prefix T404/softfloat/propagateFloat64NaN/7.3

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsp18SPILL10 for prefix T404/softfloat/propagateFloat64NaN/18.2/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tspr18.2 for prefix T404/softfloat/propagateFloat64NaN/18.2

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsp19_SPILL for prefix T404/softfloat/packFloat64/19.7/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tss23_SPILL for prefix T404/softfloat/shift64RightJamming/23.6/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tssh23.6 for prefix T404/softfloat/shift64RightJamming/23.6

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsp27SPILL10 for prefix T404/softfloat/propagateFloat64NaN/27.2/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tspr27.2 for prefix T404/softfloat/propagateFloat64NaN/27.2

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tss32_SPILL for prefix T404/softfloat/shift64RightJamming/32.5/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tssh32.5 for prefix T404/softfloat/shift64RightJamming/32.5

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsno34.9 for prefix T404/softfloat/normalizeRoundAndPackFloat64/34.9

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsr0._SPILL for prefix T404/softfloat/roundAndPackFloat64/0.16/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsro0.16 for prefix T404/softfloat/roundAndPackFloat64/0.16

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsf0SPILL14 for prefix T404/softfloat/float64_le/0.3/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tsfl0.3 for prefix T404/softfloat/float64_le/0.3

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tse5._SPILL for prefix T404/softfloat/extractFloat64Sign/5.2/_SPILL

//----------------------------------------------------------

//Report from Abbreviation:::
//Setting up abbreviation Tse5SPILL10 for prefix T404/softfloat/extractFloat64Sign/5.5/_SPILL

//----------------------------------------------------------

//Report from KiwiC-fe.rpt:::
//KiwiC: front end input processing of class or method called KiwiSystem/Kiwi
//
//root_walk start thread at a static method (used as an entry point). Method name=.cctor uid=cctor10
//
//KiwiC start_thread (or entry point) id=cctor10
//
//Root method elaborated: specificf=S_kickoff_collate leftover=1+0
//
//KiwiC: front end input processing of class or method called System/BitConverter
//
//root_walk start thread at a static method (used as an entry point). Method name=.cctor uid=cctor12
//
//KiwiC start_thread (or entry point) id=cctor12
//
//Root method elaborated: specificf=S_kickoff_collate leftover=1+1
//
//KiwiC: front end input processing of class or method called softfloat
//
//root_walk start thread at a static method (used as an entry point). Method name=.cctor uid=cctor14
//
//KiwiC start_thread (or entry point) id=cctor14
//
//Root method elaborated: specificf=S_kickoff_collate leftover=1+2
//
//KiwiC: front end input processing of class or method called dfsin
//
//root_walk start thread at a static method (used as an entry point). Method name=.cctor uid=cctor16
//
//KiwiC start_thread (or entry point) id=cctor16
//
//Root method elaborated: specificf=S_kickoff_collate leftover=1+3
//
//KiwiC: front end input processing of class or method called dfsin
//
//root_compiler: start elaborating class 'dfsin'
//
//elaborating class 'dfsin'
//
//compiling static method as entry point: style=Root idl=dfsin/Main
//
//Performing root elaboration of method Main
//
//KiwiC start_thread (or entry point) id=Main10
//
//root_compiler class done: dfsin
//
//Report of all settings used from the recipe or command line:
//
//   cil-uwind-budget=10000
//
//   kiwic-finish=enable
//
//   kiwic-cil-dump=combined
//
//   kiwic-kcode-dump=enable
//
//   kiwic-register-colours=disable
//
//   array-4d-name=KIWIARRAY4D
//
//   array-3d-name=KIWIARRAY3D
//
//   array-2d-name=KIWIARRAY2D
//
//   kiwi-dll=Kiwi.dll
//
//   kiwic-dll=Kiwic.dll
//
//   kiwic-zerolength-arrays=disable
//
//   kiwic-fpgaconsole-default=enable
//
//   postgen-optimise=enable
//
//   gtrace-loglevel=20
//
//   firstpass-loglevel=20
//
//   root=$attributeroot
//
//   ?>?=srcfile, dfsin.exe, ../softfloat.dll
//
//END OF KIWIC REPORT FILE
//

//----------------------------------------------------------

//Report from enumbers:::
//Concise expression alias report.
//
//  -- No expression aliases to report
//

//----------------------------------------------------------

//Report from verilog_render:::
//1 vectors of width 13
//
//261 vectors of width 64
//
//52 vectors of width 1
//
//30 vectors of width 16
//
//16 vectors of width 32
//
//3 vectors of width 8
//
//72 array locations of width 64
//
//259 array locations of width 8
//
//1024 bits in scalar variables
//
//Total state bits in module = 25489 bits.
//
//Total number of leaf cells = 0
//

//Major Statistics Report:
//Thread .cctor uid=cctor10 has 3 CIL instructions in 1 basic blocks
//Thread .cctor uid=cctor12 has 2 CIL instructions in 1 basic blocks
//Thread .cctor uid=cctor14 has 6 CIL instructions in 1 basic blocks
//Thread .cctor uid=cctor16 has 14 CIL instructions in 1 basic blocks
//Thread Main uid=Main10 has 2607 CIL instructions in 1010 basic blocks
//Thread mpc10 has 4930 bevelab control states (pauses)
// eof (HPR L/S Verilog)
