

// CBG Orangepath HPR L/S System

// Verilog output file generated at 22/06/2016 08:27:30
// Kiwi Scientific Acceleration (KiwiC .net/CIL/C# to Verilog/SystemC compiler): Version alpha 2.15f : 19th-June-2016 Unix 3.19.8.100
//  /home/djg11/d320/hprls/kiwipro/kiwic/distro/lib/kiwic.exe -give-backtrace -vnl=cuckoo_hash_demo.v cuckoo_hash_demo.exe -vnl-resets=synchronous -kiwic-cil-dump=combined -kiwic-kcode-dump=enable -res2-loadstore-port-count=0 -vnl-roundtrip=disable -bevelab-default-pause-mode=soft -bevelab-soft-pause-threshold=10 -vnl-rootmodname=DUT
`timescale 1ns/1ns


module DUT(output reg [639:0] KppWaypoint0, output [639:0] KppWaypoint1, output reg done, input clk, input reset);
  integer TTMT4Main_V_2;
  integer TTMT4Main_V_3;
  integer TTMT4Main_V_4;
  integer TTMT4Main_V_5;
  reg [63:0] TTMT4Main_V_6;
  integer TTMT4Main_V_7;
  integer TTMT4Main_V_8;
  integer TTMT4Main_V_9;
  integer TTMT4Main_V_10;
  integer TTMT4Main_V_11;
  reg [63:0] TTMT4Main_V_12;
  reg [63:0] TTMT4Main_V_13;
  integer TTMT4Main_V_14;
  integer TCCl0_12_V_0;
  integer TCCl0_12_V_1;
  reg [63:0] TDGe1_4_V_0;
  integer TCin1_9_V_0;
  integer TCin1_9_V_1;
  integer TCin1_9_V_2;
  integer TCin1_9_V_3;
  integer TCin1_9_V_4;
  integer TCin1_9_V_5;
  integer TCin1_9_V_6;
  integer TCin1_9_V_7;
  integer TCha6_10_V_0;
  reg [63:0] TDGe6_4_V_0;
  integer TClo6_9_V_0;
  integer TClo6_9_V_1;
  integer TClo6_9_V_2;
  integer TCha3_10_V_0;
  reg [63:0] fastspilldup30;
  integer TCl6_SPILL_256;
  reg [63:0] fastspilldup12;
  integer TCi1_SPILL_256;
  integer fastspilldup16;
  integer fastspilldup26;
  reg [63:0] A_64_US_CC_SCALbx28_dk;
  reg signed [31:0] A_sA_SINT_CC_SCALbx22_ARB0[3:0];
  reg signed [31:0] A_sA_SINT_CC_SCALbx20_ARA0[3:0];
  reg signed [31:0] A_SINT_CC_SCALbx28_seed;
  reg signed [31:0] A_SINT_CC_SCALbx24_waycap;
  reg signed [31:0] A_SINT_CC_SCALbx24_stats_lookups;
  reg signed [31:0] A_SINT_CC_SCALbx24_stats_lookup_probes;
  reg signed [31:0] A_SINT_CC_SCALbx24_next_free;
  reg signed [31:0] A_SINT_CC_SCALbx24_stats_inserts;
  reg signed [31:0] A_SINT_CC_SCALbx24_stats_insert_probes;
  reg signed [31:0] A_SINT_CC_SCALbx24_stats_insert_evictions;
  reg signed [31:0] A_SINT_CC_SCALbx24_next_victim;
  wire signed [31:0] A_SINT_CC_MAPR10NoCE3_ARA0_RDD0;
  reg [12:0] A_SINT_CC_MAPR10NoCE3_ARA0_AD0;
  reg A_SINT_CC_MAPR10NoCE3_ARA0_WEN0;
  reg A_SINT_CC_MAPR10NoCE3_ARA0_REN0;
  reg signed [31:0] A_SINT_CC_MAPR10NoCE3_ARA0_WRD0;
  wire signed [31:0] A_SINT_CC_MAPR10NoCE2_ARA0_RDD0;
  reg [12:0] A_SINT_CC_MAPR10NoCE2_ARA0_AD0;
  reg A_SINT_CC_MAPR10NoCE2_ARA0_WEN0;
  reg A_SINT_CC_MAPR10NoCE2_ARA0_REN0;
  reg signed [31:0] A_SINT_CC_MAPR10NoCE2_ARA0_WRD0;
  wire signed [31:0] A_SINT_CC_MAPR10NoCE1_ARA0_RDD0;
  reg [12:0] A_SINT_CC_MAPR10NoCE1_ARA0_AD0;
  reg A_SINT_CC_MAPR10NoCE1_ARA0_WEN0;
  reg A_SINT_CC_MAPR10NoCE1_ARA0_REN0;
  reg signed [31:0] A_SINT_CC_MAPR10NoCE1_ARA0_WRD0;
  wire signed [31:0] A_SINT_CC_MAPR10NoCE0_ARA0_RDD0;
  reg [12:0] A_SINT_CC_MAPR10NoCE0_ARA0_AD0;
  reg A_SINT_CC_MAPR10NoCE0_ARA0_WEN0;
  reg A_SINT_CC_MAPR10NoCE0_ARA0_REN0;
  reg signed [31:0] A_SINT_CC_MAPR10NoCE0_ARA0_WRD0;
  wire isMODULUS10_rdy;
  reg isMODULUS10_req;
  wire [31:0] isMODULUS10_RR;
  reg [31:0] isMODULUS10_NN;
  reg [31:0] isMODULUS10_DD;
  wire isMODULUS10_err;
  wire signed [31:0] A_SINT_CC_MAPR12NoCE3_ARB0_RDD0;
  reg [12:0] A_SINT_CC_MAPR12NoCE3_ARB0_AD0;
  reg A_SINT_CC_MAPR12NoCE3_ARB0_WEN0;
  reg A_SINT_CC_MAPR12NoCE3_ARB0_REN0;
  reg signed [31:0] A_SINT_CC_MAPR12NoCE3_ARB0_WRD0;
  wire signed [31:0] A_SINT_CC_MAPR12NoCE2_ARB0_RDD0;
  reg [12:0] A_SINT_CC_MAPR12NoCE2_ARB0_AD0;
  reg A_SINT_CC_MAPR12NoCE2_ARB0_WEN0;
  reg A_SINT_CC_MAPR12NoCE2_ARB0_REN0;
  reg signed [31:0] A_SINT_CC_MAPR12NoCE2_ARB0_WRD0;
  wire signed [31:0] A_SINT_CC_MAPR12NoCE1_ARB0_RDD0;
  reg [12:0] A_SINT_CC_MAPR12NoCE1_ARB0_AD0;
  reg A_SINT_CC_MAPR12NoCE1_ARB0_WEN0;
  reg A_SINT_CC_MAPR12NoCE1_ARB0_REN0;
  reg signed [31:0] A_SINT_CC_MAPR12NoCE1_ARB0_WRD0;
  wire signed [31:0] A_SINT_CC_MAPR12NoCE0_ARB0_RDD0;
  reg [12:0] A_SINT_CC_MAPR12NoCE0_ARB0_AD0;
  reg A_SINT_CC_MAPR12NoCE0_ARB0_WEN0;
  reg A_SINT_CC_MAPR12NoCE0_ARB0_REN0;
  reg signed [31:0] A_SINT_CC_MAPR12NoCE0_ARB0_WRD0;
  wire [63:0] A_64_US_CC_SCALbx26_ARA0_RDD0;
  reg [14:0] A_64_US_CC_SCALbx26_ARA0_AD0;
  reg A_64_US_CC_SCALbx26_ARA0_WEN0;
  reg A_64_US_CC_SCALbx26_ARA0_REN0;
  reg [63:0] A_64_US_CC_SCALbx26_ARA0_WRD0;
  reg xpc10_trk64;
  reg xpc10_trk63;
  reg xpc10_trk62;
  reg xpc10_trk61;
  reg xpc10_trk60;
  reg xpc10_trk59;
  reg xpc10_trk58;
  reg xpc10_trk57;
  reg xpc10_trk56;
  reg xpc10_trk55;
  reg xpc10_trk54;
  reg xpc10_trk53;
  reg xpc10_trk52;
  reg xpc10_trk51;
  reg xpc10_trk50;
  reg xpc10_trk49;
  reg xpc10_trk48;
  reg xpc10_trk47;
  reg xpc10_trk46;
  reg xpc10_trk45;
  reg xpc10_trk44;
  reg xpc10_trk43;
  reg xpc10_trk42;
  reg xpc10_trk41;
  reg xpc10_trk40;
  reg xpc10_trk39;
  reg xpc10_trk38;
  reg xpc10_trk37;
  reg xpc10_trk36;
  reg xpc10_trk35;
  reg xpc10_trk34;
  reg xpc10_trk33;
  reg xpc10_trk32;
  reg xpc10_trk31;
  reg xpc10_trk30;
  reg xpc10_trk29;
  reg xpc10_trk28;
  reg xpc10_trk27;
  reg xpc10_trk26;
  reg xpc10_trk25;
  reg xpc10_trk24;
  reg xpc10_trk23;
  reg xpc10_trk22;
  reg xpc10_trk21;
  reg xpc10_trk20;
  reg xpc10_trk19;
  reg xpc10_trk18;
  reg xpc10_trk17;
  reg xpc10_trk16;
  reg xpc10_trk15;
  reg xpc10_trk14;
  reg xpc10_trk13;
  reg xpc10_trk12;
  reg xpc10_trk11;
  reg xpc10_trk10;
  reg xpc10_trk9;
  reg xpc10_trk8;
  reg xpc10_trk7;
  reg xpc10_trk6;
  reg xpc10_trk5;
  reg xpc10_trk4;
  reg xpc10_trk3;
  reg xpc10_trk2;
  reg xpc10_trk1;
  reg xpc10_trk0;
  reg xpc10_stall;
  reg xpc10_clear;
  reg [63:0] Z64USCCSCALbx26ARA0RRh10hold;
  reg Z64USCCSCALbx26ARA0RRh10shot0;
  reg signed [31:0] SINTCCMAPR12NoCE0ARB0RRh10hold;
  reg SINTCCMAPR12NoCE0ARB0RRh10shot0;
  reg signed [31:0] SINTCCMAPR12NoCE1ARB0RRh10hold;
  reg SINTCCMAPR12NoCE1ARB0RRh10shot0;
  reg signed [31:0] SINTCCMAPR12NoCE2ARB0RRh10hold;
  reg SINTCCMAPR12NoCE2ARB0RRh10shot0;
  reg signed [31:0] SINTCCMAPR12NoCE3ARB0RRh10hold;
  reg SINTCCMAPR12NoCE3ARB0RRh10shot0;
  reg signed [31:0] SINTCCMAPR10NoCE0ARA0RRh10hold;
  reg SINTCCMAPR10NoCE0ARA0RRh10shot0;
  reg signed [31:0] SINTCCMAPR10NoCE1ARA0RRh10hold;
  reg SINTCCMAPR10NoCE1ARA0RRh10shot0;
  reg signed [31:0] SINTCCMAPR10NoCE2ARA0RRh10hold;
  reg SINTCCMAPR10NoCE2ARA0RRh10shot0;
  reg signed [31:0] SINTCCMAPR10NoCE3ARA0RRh10hold;
  reg SINTCCMAPR10NoCE3ARA0RRh10shot0;
  reg isMODULUS10RRh10primed;
  reg isMODULUS10RRh10vld;
  reg signed [31:0] isMODULUS10RRh10hold;
  reg [9:0] xpc10nz;
 always   @(* )  begin 
       KppWaypoint0 = 0;
       A_SINT_CC_MAPR12NoCE3_ARB0_WRD0 = 0;
       A_SINT_CC_MAPR12NoCE2_ARB0_WRD0 = 0;
       A_SINT_CC_MAPR12NoCE1_ARB0_WRD0 = 0;
       A_SINT_CC_MAPR12NoCE0_ARB0_WRD0 = 0;
       A_64_US_CC_SCALbx26_ARA0_WRD0 = 0;
       A_64_US_CC_SCALbx26_ARA0_AD0 = 0;
       A_SINT_CC_MAPR12NoCE0_ARB0_AD0 = 0;
       A_SINT_CC_MAPR12NoCE1_ARB0_AD0 = 0;
       A_SINT_CC_MAPR12NoCE2_ARB0_AD0 = 0;
       A_SINT_CC_MAPR12NoCE3_ARB0_AD0 = 0;
       isMODULUS10_NN = 0;
       isMODULUS10_DD = 0;
       A_SINT_CC_MAPR10NoCE3_ARA0_AD0 = 0;
       A_SINT_CC_MAPR10NoCE3_ARA0_WRD0 = 0;
       A_SINT_CC_MAPR10NoCE2_ARA0_AD0 = 0;
       A_SINT_CC_MAPR10NoCE2_ARA0_WRD0 = 0;
       A_SINT_CC_MAPR10NoCE1_ARA0_AD0 = 0;
       A_SINT_CC_MAPR10NoCE1_ARA0_WRD0 = 0;
       A_SINT_CC_MAPR10NoCE0_ARA0_AD0 = 0;
       A_SINT_CC_MAPR10NoCE0_ARA0_WRD0 = 0;
       A_SINT_CC_MAPR10NoCE3_ARA0_WEN0 = 0;
       A_SINT_CC_MAPR10NoCE2_ARA0_WEN0 = 0;
       A_SINT_CC_MAPR10NoCE1_ARA0_WEN0 = 0;
       A_SINT_CC_MAPR10NoCE0_ARA0_WEN0 = 0;
       A_SINT_CC_MAPR12NoCE3_ARB0_WEN0 = 0;
       A_SINT_CC_MAPR12NoCE2_ARB0_WEN0 = 0;
       A_SINT_CC_MAPR12NoCE1_ARB0_WEN0 = 0;
       A_SINT_CC_MAPR12NoCE0_ARB0_WEN0 = 0;
       A_SINT_CC_MAPR10NoCE0_ARA0_REN0 = 0;
       A_SINT_CC_MAPR10NoCE1_ARA0_REN0 = 0;
       A_SINT_CC_MAPR10NoCE2_ARA0_REN0 = 0;
       A_SINT_CC_MAPR10NoCE3_ARA0_REN0 = 0;
       isMODULUS10_req = 0;
       A_SINT_CC_MAPR12NoCE0_ARB0_REN0 = 0;
       A_SINT_CC_MAPR12NoCE1_ARB0_REN0 = 0;
       A_SINT_CC_MAPR12NoCE2_ARB0_REN0 = 0;
       A_SINT_CC_MAPR12NoCE3_ARB0_REN0 = 0;
       A_64_US_CC_SCALbx26_ARA0_WEN0 = 0;
       A_64_US_CC_SCALbx26_ARA0_REN0 = 0;
      if (!xpc10_stall)  begin 
               A_64_US_CC_SCALbx26_ARA0_REN0 = ((xpc10nz==8'd239/*US*/)? 1'd1: 1'd0);
               A_64_US_CC_SCALbx26_ARA0_WEN0 = ((xpc10nz==8'd255/*US*/)? 1'd1: 1'd0);
               A_SINT_CC_MAPR12NoCE3_ARB0_REN0 = ((xpc10nz==8'd236/*US*/) && (TTMT4Main_V_11==((A_sA_SINT_CC_SCALbx20_ARA0[TClo6_9_V_0
              ]==2'd3/*MS*/)? ((xpc10nz==8'd237/*US*/)? A_SINT_CC_MAPR10NoCE3_ARA0_RDD0: SINTCCMAPR10NoCE3ARA0RRh10hold): ((A_sA_SINT_CC_SCALbx20_ARA0
              [TClo6_9_V_0]==2'd2/*MS*/)? ((xpc10nz==8'd237/*US*/)? A_SINT_CC_MAPR10NoCE2_ARA0_RDD0: SINTCCMAPR10NoCE2ARA0RRh10hold): ((A_sA_SINT_CC_SCALbx20_ARA0
              [TClo6_9_V_0]==1'd1/*MS*/)? ((xpc10nz==8'd237/*US*/)? A_SINT_CC_MAPR10NoCE1_ARA0_RDD0: SINTCCMAPR10NoCE1ARA0RRh10hold): ((A_sA_SINT_CC_SCALbx20_ARA0
              [TClo6_9_V_0]==0/*MS*/)? ((xpc10nz==8'd237/*US*/)? A_SINT_CC_MAPR10NoCE0_ARA0_RDD0: SINTCCMAPR10NoCE0ARA0RRh10hold): 1'bx
              ))))) || (TClo6_9_V_0>=3'd4) && (xpc10nz==8'd242/*US*/)) && (TClo6_9_V_0!=3'd4/*US*/) || (xpc10nz==9'd287/*US*/);

               A_SINT_CC_MAPR12NoCE2_ARB0_REN0 = ((xpc10nz==8'd236/*US*/) && (TTMT4Main_V_11==((A_sA_SINT_CC_SCALbx20_ARA0[TClo6_9_V_0
              ]==2'd3/*MS*/)? ((xpc10nz==8'd237/*US*/)? A_SINT_CC_MAPR10NoCE3_ARA0_RDD0: SINTCCMAPR10NoCE3ARA0RRh10hold): ((A_sA_SINT_CC_SCALbx20_ARA0
              [TClo6_9_V_0]==2'd2/*MS*/)? ((xpc10nz==8'd237/*US*/)? A_SINT_CC_MAPR10NoCE2_ARA0_RDD0: SINTCCMAPR10NoCE2ARA0RRh10hold): ((A_sA_SINT_CC_SCALbx20_ARA0
              [TClo6_9_V_0]==1'd1/*MS*/)? ((xpc10nz==8'd237/*US*/)? A_SINT_CC_MAPR10NoCE1_ARA0_RDD0: SINTCCMAPR10NoCE1ARA0RRh10hold): ((A_sA_SINT_CC_SCALbx20_ARA0
              [TClo6_9_V_0]==0/*MS*/)? ((xpc10nz==8'd237/*US*/)? A_SINT_CC_MAPR10NoCE0_ARA0_RDD0: SINTCCMAPR10NoCE0ARA0RRh10hold): 1'bx
              ))))) || (TClo6_9_V_0>=3'd4) && (xpc10nz==8'd242/*US*/)) && (TClo6_9_V_0!=3'd4/*US*/) || (xpc10nz==9'd287/*US*/);

               A_SINT_CC_MAPR12NoCE1_ARB0_REN0 = ((xpc10nz==8'd236/*US*/) && (TTMT4Main_V_11==((A_sA_SINT_CC_SCALbx20_ARA0[TClo6_9_V_0
              ]==2'd3/*MS*/)? ((xpc10nz==8'd237/*US*/)? A_SINT_CC_MAPR10NoCE3_ARA0_RDD0: SINTCCMAPR10NoCE3ARA0RRh10hold): ((A_sA_SINT_CC_SCALbx20_ARA0
              [TClo6_9_V_0]==2'd2/*MS*/)? ((xpc10nz==8'd237/*US*/)? A_SINT_CC_MAPR10NoCE2_ARA0_RDD0: SINTCCMAPR10NoCE2ARA0RRh10hold): ((A_sA_SINT_CC_SCALbx20_ARA0
              [TClo6_9_V_0]==1'd1/*MS*/)? ((xpc10nz==8'd237/*US*/)? A_SINT_CC_MAPR10NoCE1_ARA0_RDD0: SINTCCMAPR10NoCE1ARA0RRh10hold): ((A_sA_SINT_CC_SCALbx20_ARA0
              [TClo6_9_V_0]==0/*MS*/)? ((xpc10nz==8'd237/*US*/)? A_SINT_CC_MAPR10NoCE0_ARA0_RDD0: SINTCCMAPR10NoCE0ARA0RRh10hold): 1'bx
              ))))) || (TClo6_9_V_0>=3'd4) && (xpc10nz==8'd242/*US*/)) && (TClo6_9_V_0!=3'd4/*US*/) || (xpc10nz==9'd287/*US*/);

               A_SINT_CC_MAPR12NoCE0_ARB0_REN0 = ((xpc10nz==8'd236/*US*/) && (TTMT4Main_V_11==((A_sA_SINT_CC_SCALbx20_ARA0[TClo6_9_V_0
              ]==2'd3/*MS*/)? ((xpc10nz==8'd237/*US*/)? A_SINT_CC_MAPR10NoCE3_ARA0_RDD0: SINTCCMAPR10NoCE3ARA0RRh10hold): ((A_sA_SINT_CC_SCALbx20_ARA0
              [TClo6_9_V_0]==2'd2/*MS*/)? ((xpc10nz==8'd237/*US*/)? A_SINT_CC_MAPR10NoCE2_ARA0_RDD0: SINTCCMAPR10NoCE2ARA0RRh10hold): ((A_sA_SINT_CC_SCALbx20_ARA0
              [TClo6_9_V_0]==1'd1/*MS*/)? ((xpc10nz==8'd237/*US*/)? A_SINT_CC_MAPR10NoCE1_ARA0_RDD0: SINTCCMAPR10NoCE1ARA0RRh10hold): ((A_sA_SINT_CC_SCALbx20_ARA0
              [TClo6_9_V_0]==0/*MS*/)? ((xpc10nz==8'd237/*US*/)? A_SINT_CC_MAPR10NoCE0_ARA0_RDD0: SINTCCMAPR10NoCE0ARA0RRh10hold): 1'bx
              ))))) || (TClo6_9_V_0>=3'd4) && (xpc10nz==8'd242/*US*/)) && (TClo6_9_V_0!=3'd4/*US*/) || (xpc10nz==9'd287/*US*/);

               isMODULUS10_req = ((TCha6_10_V_0>=0) && (xpc10nz==9'd342/*US*/) || (TCha3_10_V_0>=0) && (xpc10nz==7'd106/*US*/) || (xpc10nz
              ==8'd171/*US*/) || (xpc10nz==9'd407/*US*/)? 1'd1: 1'd0);

               A_SINT_CC_MAPR10NoCE3_ARA0_REN0 = ((xpc10nz==9'd285/*US*/) || (xpc10nz==8'd236/*US*/) || (xpc10nz==9'd472/*US*/)? 1'd1
              : 1'd0);

               A_SINT_CC_MAPR10NoCE2_ARA0_REN0 = ((xpc10nz==9'd285/*US*/) || (xpc10nz==8'd236/*US*/) || (xpc10nz==9'd472/*US*/)? 1'd1
              : 1'd0);

               A_SINT_CC_MAPR10NoCE1_ARA0_REN0 = ((xpc10nz==9'd285/*US*/) || (xpc10nz==8'd236/*US*/) || (xpc10nz==9'd472/*US*/)? 1'd1
              : 1'd0);

               A_SINT_CC_MAPR10NoCE0_ARA0_REN0 = ((xpc10nz==9'd285/*US*/) || (xpc10nz==8'd236/*US*/) || (xpc10nz==9'd472/*US*/)? 1'd1
              : 1'd0);

               A_SINT_CC_MAPR12NoCE0_ARB0_WEN0 = ((xpc10nz==9'd327/*US*/) || (xpc10nz==9'd314/*US*/) || (xpc10nz==9'd324/*US*/) || (((A_sA_SINT_CC_SCALbx20_ARA0
              [A_SINT_CC_SCALbx24_next_victim]==2'd3/*MS*/)? 1'd1: (A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]!=0/*MS*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim
              ]!=2'd2/*MS*/)) || (A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]==0/*MS*/) || (A_sA_SINT_CC_SCALbx20_ARA0
              [A_SINT_CC_SCALbx24_next_victim]==1'd1/*MS*/) || (A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]==2'd2/*MS*/)) && 
              (xpc10nz==9'd289/*US*/)) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]==0/*MS*/) || (((((A_sA_SINT_CC_SCALbx20_ARA0
              [TCin1_9_V_4]==2'd3/*MS*/)? (xpc10nz==9'd503/*US*/) || (xpc10nz==9'd259/*US*/): ((xpc10nz==9'd503/*US*/) || (xpc10nz==9'd259
              /*US*/)) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=1'd1/*MS*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd2/*MS*/)) || ((xpc10nz==9'd503/*US*/) || (xpc10nz==9'd259/*US*/)) && (A_sA_SINT_CC_SCALbx20_ARA0
              [TCin1_9_V_4]==0/*MS*/) || ((xpc10nz==9'd503/*US*/) || (xpc10nz==9'd259/*US*/)) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4
              ]==1'd1/*MS*/) || ((xpc10nz==9'd503/*US*/) || (xpc10nz==9'd259/*US*/)) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd2
              /*MS*/)) && (TCin1_9_V_4>=3'd4) || ((A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd3/*MS*/)? !A_SINT_CC_MAPR10NoCE3_ARA0_RDD0
               && (xpc10nz==9'd473/*US*/): (xpc10nz==9'd473/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd2/*MS*/)) || !A_SINT_CC_MAPR10NoCE0_ARA0_RDD0
               && (xpc10nz==9'd473/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==0/*MS*/) || !A_SINT_CC_MAPR10NoCE1_ARA0_RDD0 && 
              (xpc10nz==9'd473/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==1'd1/*MS*/) || !A_SINT_CC_MAPR10NoCE2_ARA0_RDD0 && 
              (xpc10nz==9'd473/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd2/*MS*/)) && (TCin1_9_V_4!=3'd4/*US*/) || (xpc10nz
              ==9'd335/*US*/) || (xpc10nz==9'd330/*US*/) || (xpc10nz==9'd338/*US*/)) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==0/*MS*/);

               A_SINT_CC_MAPR12NoCE1_ARB0_WEN0 = ((xpc10nz==9'd314/*US*/) || (xpc10nz==9'd324/*US*/) || (((A_sA_SINT_CC_SCALbx20_ARA0
              [A_SINT_CC_SCALbx24_next_victim]==2'd3/*MS*/)? 1'd1: (A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]!=0/*MS*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim
              ]!=2'd2/*MS*/)) || (A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]==0/*MS*/) || (A_sA_SINT_CC_SCALbx20_ARA0
              [A_SINT_CC_SCALbx24_next_victim]==1'd1/*MS*/) || (A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]==2'd2/*MS*/)) && 
              (xpc10nz==9'd289/*US*/)) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]==1'd1/*MS*/) || (((((A_sA_SINT_CC_SCALbx20_ARA0
              [TCin1_9_V_4]==2'd3/*MS*/)? (xpc10nz==9'd503/*US*/) || (xpc10nz==9'd259/*US*/): ((xpc10nz==9'd503/*US*/) || (xpc10nz==9'd259
              /*US*/)) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=1'd1/*MS*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd2/*MS*/)) || ((xpc10nz==9'd503/*US*/) || (xpc10nz==9'd259/*US*/)) && (A_sA_SINT_CC_SCALbx20_ARA0
              [TCin1_9_V_4]==0/*MS*/) || ((xpc10nz==9'd503/*US*/) || (xpc10nz==9'd259/*US*/)) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4
              ]==1'd1/*MS*/) || ((xpc10nz==9'd503/*US*/) || (xpc10nz==9'd259/*US*/)) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd2
              /*MS*/)) && (TCin1_9_V_4>=3'd4) || ((A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd3/*MS*/)? !A_SINT_CC_MAPR10NoCE3_ARA0_RDD0
               && (xpc10nz==9'd473/*US*/): (xpc10nz==9'd473/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd2/*MS*/)) || !A_SINT_CC_MAPR10NoCE0_ARA0_RDD0
               && (xpc10nz==9'd473/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==0/*MS*/) || !A_SINT_CC_MAPR10NoCE1_ARA0_RDD0 && 
              (xpc10nz==9'd473/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==1'd1/*MS*/) || !A_SINT_CC_MAPR10NoCE2_ARA0_RDD0 && 
              (xpc10nz==9'd473/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd2/*MS*/)) && (TCin1_9_V_4!=3'd4/*US*/) || (xpc10nz
              ==9'd330/*US*/) || (xpc10nz==9'd335/*US*/)) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==1'd1/*MS*/);

               A_SINT_CC_MAPR12NoCE2_ARB0_WEN0 = ((xpc10nz==9'd314/*US*/) || (((A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim
              ]==2'd3/*MS*/)? 1'd1: (A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [A_SINT_CC_SCALbx24_next_victim]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]!=2'd2/*MS*/)) || 
              (A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]==0/*MS*/) || (A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim
              ]==1'd1/*MS*/) || (A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]==2'd2/*MS*/)) && (xpc10nz==9'd289/*US*/)) && 
              (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]==2'd2/*MS*/) || (((((A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4
              ]==2'd3/*MS*/)? (xpc10nz==9'd503/*US*/) || (xpc10nz==9'd259/*US*/): ((xpc10nz==9'd503/*US*/) || (xpc10nz==9'd259/*US*/)) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [TCin1_9_V_4]!=2'd2/*MS*/)) || ((xpc10nz==9'd503/*US*/) || (xpc10nz==9'd259/*US*/)) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4
              ]==0/*MS*/) || ((xpc10nz==9'd503/*US*/) || (xpc10nz==9'd259/*US*/)) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==1'd1/*MS*/) || 
              ((xpc10nz==9'd503/*US*/) || (xpc10nz==9'd259/*US*/)) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd2/*MS*/)) && (TCin1_9_V_4
              >=3'd4) || ((A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd3/*MS*/)? !A_SINT_CC_MAPR10NoCE3_ARA0_RDD0 && (xpc10nz==9'd473
              /*US*/): (xpc10nz==9'd473/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4
              ]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd2/*MS*/)) || !A_SINT_CC_MAPR10NoCE0_ARA0_RDD0 && (xpc10nz
              ==9'd473/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==0/*MS*/) || !A_SINT_CC_MAPR10NoCE1_ARA0_RDD0 && (xpc10nz==
              9'd473/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==1'd1/*MS*/) || !A_SINT_CC_MAPR10NoCE2_ARA0_RDD0 && (xpc10nz==
              9'd473/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd2/*MS*/)) && (TCin1_9_V_4!=3'd4/*US*/) || (xpc10nz==9'd330
              /*US*/)) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd2/*MS*/);

               A_SINT_CC_MAPR12NoCE3_ARB0_WEN0 = ((((A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd3/*MS*/)? (xpc10nz==9'd503/*US*/) || 
              (xpc10nz==9'd259/*US*/): ((xpc10nz==9'd503/*US*/) || (xpc10nz==9'd259/*US*/)) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4
              ]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd2/*MS*/)) || 
              ((xpc10nz==9'd503/*US*/) || (xpc10nz==9'd259/*US*/)) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==0/*MS*/) || ((xpc10nz
              ==9'd503/*US*/) || (xpc10nz==9'd259/*US*/)) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==1'd1/*MS*/) || ((xpc10nz==9'd503
              /*US*/) || (xpc10nz==9'd259/*US*/)) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd2/*MS*/)) && (TCin1_9_V_4>=3'd4) || 
              ((A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd3/*MS*/)? !A_SINT_CC_MAPR10NoCE3_ARA0_RDD0 && (xpc10nz==9'd473/*US*/): (xpc10nz
              ==9'd473/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=1'd1
              /*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd2/*MS*/)) || !A_SINT_CC_MAPR10NoCE0_ARA0_RDD0 && (xpc10nz==9'd473
              /*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==0/*MS*/) || !A_SINT_CC_MAPR10NoCE1_ARA0_RDD0 && (xpc10nz==9'd473/*US*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==1'd1/*MS*/) || !A_SINT_CC_MAPR10NoCE2_ARA0_RDD0 && (xpc10nz==9'd473/*US*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd2/*MS*/)) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd3/*MS*/) && (TCin1_9_V_4
              !=3'd4/*US*/) || (((A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]==2'd3/*MS*/)? 1'd1: (A_sA_SINT_CC_SCALbx20_ARA0
              [A_SINT_CC_SCALbx24_next_victim]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]!=1'd1/*MS*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]!=2'd2/*MS*/)) || (A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim
              ]==0/*MS*/) || (A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]==1'd1/*MS*/) || (A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim
              ]==2'd2/*MS*/)) && (xpc10nz==9'd289/*US*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]==2'd3/*MS*/);

               A_SINT_CC_MAPR10NoCE0_ARA0_WEN0 = ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==0/*MS*/)? (((xpc10nz==5'd20/*US*/) || (xpc10nz==
              7'd65/*US*/) && (TCCl0_12_V_0<A_SINT_CC_SCALbx24_waycap)) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) || ((xpc10nz==6'd37/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [1'd1]!=2'd3/*MS*/) || (xpc10nz==10'd576/*US*/)) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) || (xpc10nz==10'd588
              /*US*/)) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) || (xpc10nz==
              10'd609/*US*/) || (xpc10nz==6'd50/*US*/) || (xpc10nz==10'd599/*US*/) || (xpc10nz==10'd550/*US*/) || (xpc10nz==10'd558/*US*/) || 
              (xpc10nz==10'd565/*US*/): (((((xpc10nz==5'd20/*US*/) || (xpc10nz==7'd65/*US*/) && (TCCl0_12_V_0<A_SINT_CC_SCALbx24_waycap
              )) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [0]!=0/*MS*/) || ((xpc10nz==6'd37/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) || (xpc10nz==10'd576/*US*/)) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) || (xpc10nz==10'd588/*US*/)) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) || 
              (xpc10nz==10'd599/*US*/)) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) || ((xpc10nz==10'd609/*US*/) || 
              (xpc10nz==6'd50/*US*/)) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) || (xpc10nz==10'd550/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) || (xpc10nz==10'd558/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) || 
              (xpc10nz==10'd565/*US*/)) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==0/*MS*/)) || ((TCin1_9_V_4==3'd4/*US*/)? !A_SINT_CC_MAPR10NoCE0_ARA0_RDD0
               && (xpc10nz==9'd473/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==0/*MS*/): ((((A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4
              ]==2'd3/*MS*/)? (xpc10nz==9'd503/*US*/) || (xpc10nz==9'd259/*US*/): ((xpc10nz==9'd503/*US*/) || (xpc10nz==9'd259/*US*/)) && 
              (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
              [TCin1_9_V_4]!=2'd2/*MS*/)) || ((xpc10nz==9'd503/*US*/) || (xpc10nz==9'd259/*US*/)) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4
              ]==0/*MS*/) || ((xpc10nz==9'd503/*US*/) || (xpc10nz==9'd259/*US*/)) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==1'd1/*MS*/) || 
              ((xpc10nz==9'd503/*US*/) || (xpc10nz==9'd259/*US*/)) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd2/*MS*/)) && (TCin1_9_V_4
              >=3'd4) || ((A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd3/*MS*/)? !A_SINT_CC_MAPR10NoCE0_ARA0_RDD0 && (xpc10nz==9'd473
              /*US*/): !A_SINT_CC_MAPR10NoCE0_ARA0_RDD0 && (xpc10nz==9'd473/*US*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=0/*MS*/) && 
              (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd2/*MS*/)) || !A_SINT_CC_MAPR10NoCE0_ARA0_RDD0
               && (xpc10nz==9'd473/*US*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==0/*MS*/) || !A_SINT_CC_MAPR10NoCE0_ARA0_RDD0 && 
              (xpc10nz==9'd473/*US*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==1'd1/*MS*/) || !A_SINT_CC_MAPR10NoCE0_ARA0_RDD0 && 
              (xpc10nz==9'd473/*US*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd2/*MS*/)) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4
              ]==0/*MS*/)) || ((xpc10nz==10'd534/*US*/) || (xpc10nz==10'd528/*US*/) || (TCCl0_12_V_1<3'd4) && (xpc10nz==10'd532/*US*/) || 
              (xpc10nz==10'd537/*US*/)) && (A_sA_SINT_CC_SCALbx20_ARA0[TCCl0_12_V_1]==0/*MS*/) || (((A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim
              ]==2'd3/*MS*/)? 1'd1: (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
              [A_SINT_CC_SCALbx24_next_victim]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]!=2'd2/*MS*/)) || 
              (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]==0/*MS*/) || (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim
              ]==1'd1/*MS*/) || (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]==2'd2/*MS*/)) && (xpc10nz==9'd289/*US*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]==0/*MS*/) || ((xpc10nz==5'd20/*US*/) || (xpc10nz==7'd65/*US*/) && 
              (TCCl0_12_V_0<A_SINT_CC_SCALbx24_waycap)) && (A_sA_SINT_CC_SCALbx20_ARA0[0]==0/*MS*/) || (((xpc10nz==5'd20/*US*/) || (xpc10nz
              ==7'd65/*US*/) && (TCCl0_12_V_0<A_SINT_CC_SCALbx24_waycap)) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) || (xpc10nz
              ==10'd599/*US*/) || (xpc10nz==10'd588/*US*/) || (xpc10nz==10'd576/*US*/) || (xpc10nz==6'd37/*US*/)) && (A_sA_SINT_CC_SCALbx20_ARA0
              [1'd1]==0/*MS*/) || ((xpc10nz==10'd547/*US*/) || (xpc10nz==10'd540/*US*/) || (xpc10nz==6'd59/*US*/) || (xpc10nz==10'd544
              /*US*/) || (xpc10nz==10'd571/*US*/) || (xpc10nz==10'd565/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==1'd1/*MS*/) || ((xpc10nz
              ==10'd558/*US*/) || (xpc10nz==10'd565/*US*/)) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==2'd2/*MS*/) || ((xpc10nz==10'd550/*US*/) || 
              (xpc10nz==10'd558/*US*/) || (xpc10nz==10'd565/*US*/)) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==2'd3/*MS*/)) && (A_sA_SINT_CC_SCALbx20_ARA0
              [2'd3]==0/*MS*/);

               A_SINT_CC_MAPR10NoCE1_ARA0_WEN0 = ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==1'd1/*MS*/)? (((xpc10nz==5'd20/*US*/) || (xpc10nz
              ==7'd65/*US*/) && (TCCl0_12_V_0<A_SINT_CC_SCALbx24_waycap)) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=1'd1/*MS*/) || ((xpc10nz==6'd37/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [1'd1]!=2'd3/*MS*/) || (xpc10nz==10'd576/*US*/)) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) || (xpc10nz==10'd588
              /*US*/)) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) || (xpc10nz==
              10'd599/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) || (xpc10nz==10'd609/*US*/) || (xpc10nz==6'd50/*US*/) || 
              (xpc10nz==10'd550/*US*/) || (xpc10nz==10'd558/*US*/) || (xpc10nz==10'd565/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==
              1'd1/*MS*/): ((((xpc10nz==5'd20/*US*/) || (xpc10nz==7'd65/*US*/) && (TCCl0_12_V_0<A_SINT_CC_SCALbx24_waycap)) && (A_sA_SINT_CC_SCALbx20_ARA0
              [1'd1]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=1'd1/*MS*/) || ((xpc10nz
              ==6'd37/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) || (xpc10nz==10'd576/*US*/)) && (A_sA_SINT_CC_SCALbx20_ARA0
              [1'd1]!=2'd2/*MS*/) || (xpc10nz==10'd588/*US*/)) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) || (xpc10nz==10'd599/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [1'd1]!=0/*MS*/) || ((xpc10nz==10'd609/*US*/) || (xpc10nz==6'd50/*US*/)) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) || (xpc10nz==10'd550/*US*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) || (xpc10nz==10'd558/*US*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/)) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==1'd1/*MS*/)) || ((TCin1_9_V_4==3'd4/*US*/)? !A_SINT_CC_MAPR10NoCE1_ARA0_RDD0
               && (xpc10nz==9'd473/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==1'd1/*MS*/): ((((A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4
              ]==2'd3/*MS*/)? (xpc10nz==9'd503/*US*/) || (xpc10nz==9'd259/*US*/): ((xpc10nz==9'd503/*US*/) || (xpc10nz==9'd259/*US*/)) && 
              (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
              [TCin1_9_V_4]!=2'd2/*MS*/)) || ((xpc10nz==9'd503/*US*/) || (xpc10nz==9'd259/*US*/)) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4
              ]==0/*MS*/) || ((xpc10nz==9'd503/*US*/) || (xpc10nz==9'd259/*US*/)) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==1'd1/*MS*/) || 
              ((xpc10nz==9'd503/*US*/) || (xpc10nz==9'd259/*US*/)) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd2/*MS*/)) && (TCin1_9_V_4
              >=3'd4) || ((A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd3/*MS*/)? !A_SINT_CC_MAPR10NoCE1_ARA0_RDD0 && (xpc10nz==9'd473
              /*US*/): !A_SINT_CC_MAPR10NoCE1_ARA0_RDD0 && (xpc10nz==9'd473/*US*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=0/*MS*/) && 
              (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd2/*MS*/)) || !A_SINT_CC_MAPR10NoCE1_ARA0_RDD0
               && (xpc10nz==9'd473/*US*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==0/*MS*/) || !A_SINT_CC_MAPR10NoCE1_ARA0_RDD0 && 
              (xpc10nz==9'd473/*US*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==1'd1/*MS*/) || !A_SINT_CC_MAPR10NoCE1_ARA0_RDD0 && 
              (xpc10nz==9'd473/*US*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd2/*MS*/)) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4
              ]==1'd1/*MS*/)) || ((xpc10nz==10'd534/*US*/) || (xpc10nz==10'd528/*US*/) || (TCCl0_12_V_1<3'd4) && (xpc10nz==10'd532/*US*/)) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[TCCl0_12_V_1]==1'd1/*MS*/) || (((A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]
              ==2'd3/*MS*/)? 1'd1: (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
              [A_SINT_CC_SCALbx24_next_victim]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]!=2'd2/*MS*/)) || 
              (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]==0/*MS*/) || (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim
              ]==1'd1/*MS*/) || (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]==2'd2/*MS*/)) && (xpc10nz==9'd289/*US*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]==1'd1/*MS*/) || ((xpc10nz==5'd20/*US*/) || (xpc10nz==7'd65/*US*/) && 
              (TCCl0_12_V_0<A_SINT_CC_SCALbx24_waycap)) && (A_sA_SINT_CC_SCALbx20_ARA0[0]==1'd1/*MS*/) || (((xpc10nz==5'd20/*US*/) || 
              (xpc10nz==7'd65/*US*/) && (TCCl0_12_V_0<A_SINT_CC_SCALbx24_waycap)) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=1'd1/*MS*/) || (xpc10nz
              ==10'd588/*US*/) || (xpc10nz==10'd576/*US*/) || (xpc10nz==6'd37/*US*/)) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]==1'd1/*MS*/) || 
              ((xpc10nz==10'd565/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) || (xpc10nz==10'd571/*US*/) || (xpc10nz==10'd544
              /*US*/) || (xpc10nz==6'd59/*US*/) || (xpc10nz==10'd540/*US*/) || ((xpc10nz==10'd565/*US*/) || (xpc10nz==10'd558/*US*/)) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==2'd2/*MS*/) || ((xpc10nz==10'd550/*US*/) || (xpc10nz==10'd565/*US*/) || (xpc10nz==10'd558
              /*US*/)) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==2'd3/*MS*/)) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==1'd1/*MS*/);

               A_SINT_CC_MAPR10NoCE2_ARA0_WEN0 = ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==2'd2/*MS*/)? (((xpc10nz==5'd20/*US*/) || (xpc10nz
              ==7'd65/*US*/) && (TCCl0_12_V_0<A_SINT_CC_SCALbx24_waycap)) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [0]!=2'd2/*MS*/) || (xpc10nz==6'd37/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) || (xpc10nz==10'd576/*US*/)) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [1'd1]!=2'd2/*MS*/) || ((xpc10nz==10'd588/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) || (xpc10nz==10'd599
              /*US*/)) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) || (xpc10nz==10'd609/*US*/) || (xpc10nz==6'd50/*US*/) || (xpc10nz
              ==10'd550/*US*/) || ((xpc10nz==10'd558/*US*/) || (xpc10nz==10'd565/*US*/)) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==2'd2/*MS*/): ((((xpc10nz
              ==5'd20/*US*/) || (xpc10nz==7'd65/*US*/) && (TCCl0_12_V_0<A_SINT_CC_SCALbx24_waycap)) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1
              ]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) || (xpc10nz==6'd37/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [1'd1]!=2'd3/*MS*/) || (xpc10nz==10'd576/*US*/)) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) || ((xpc10nz==10'd588/*US*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) || (xpc10nz==10'd599/*US*/)) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [1'd1]!=0/*MS*/) || ((xpc10nz==10'd609/*US*/) || (xpc10nz==6'd50/*US*/)) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) || (xpc10nz==10'd550/*US*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/)) && (A_sA_SINT_CC_SCALbx20_ARA0
              [2'd3]==2'd2/*MS*/)) || ((TCin1_9_V_4==3'd4/*US*/)? !A_SINT_CC_MAPR10NoCE2_ARA0_RDD0 && (xpc10nz==9'd473/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [TCin1_9_V_4]==2'd2/*MS*/): ((((A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd3/*MS*/)? (xpc10nz==9'd503/*US*/) || (xpc10nz
              ==9'd259/*US*/): ((xpc10nz==9'd503/*US*/) || (xpc10nz==9'd259/*US*/)) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=0/*MS*/) && 
              (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd2/*MS*/)) || ((xpc10nz
              ==9'd503/*US*/) || (xpc10nz==9'd259/*US*/)) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==0/*MS*/) || ((xpc10nz==9'd503/*US*/) || 
              (xpc10nz==9'd259/*US*/)) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==1'd1/*MS*/) || ((xpc10nz==9'd503/*US*/) || (xpc10nz
              ==9'd259/*US*/)) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd2/*MS*/)) && (TCin1_9_V_4>=3'd4) || ((A_sA_SINT_CC_SCALbx22_ARB0
              [TCin1_9_V_4]==2'd3/*MS*/)? !A_SINT_CC_MAPR10NoCE2_ARA0_RDD0 && (xpc10nz==9'd473/*US*/): !A_SINT_CC_MAPR10NoCE2_ARA0_RDD0
               && (xpc10nz==9'd473/*US*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4
              ]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd2/*MS*/)) || !A_SINT_CC_MAPR10NoCE2_ARA0_RDD0 && (xpc10nz
              ==9'd473/*US*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==0/*MS*/) || !A_SINT_CC_MAPR10NoCE2_ARA0_RDD0 && (xpc10nz==
              9'd473/*US*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==1'd1/*MS*/) || !A_SINT_CC_MAPR10NoCE2_ARA0_RDD0 && (xpc10nz==
              9'd473/*US*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd2/*MS*/)) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd2
              /*MS*/)) || ((xpc10nz==10'd528/*US*/) || (TCCl0_12_V_1<3'd4) && (xpc10nz==10'd532/*US*/)) && (A_sA_SINT_CC_SCALbx20_ARA0
              [TCCl0_12_V_1]==2'd2/*MS*/) || (((A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]==2'd3/*MS*/)? 1'd1: (A_sA_SINT_CC_SCALbx22_ARB0
              [A_SINT_CC_SCALbx24_next_victim]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]!=1'd1/*MS*/) && 
              (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]!=2'd2/*MS*/)) || (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim
              ]==0/*MS*/) || (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]==1'd1/*MS*/) || (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim
              ]==2'd2/*MS*/)) && (xpc10nz==9'd289/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]==2'd2/*MS*/) || 
              ((xpc10nz==5'd20/*US*/) || (xpc10nz==7'd65/*US*/) && (TCCl0_12_V_0<A_SINT_CC_SCALbx24_waycap)) && (A_sA_SINT_CC_SCALbx20_ARA0
              [0]==2'd2/*MS*/) || (((xpc10nz==5'd20/*US*/) || (xpc10nz==7'd65/*US*/) && (TCCl0_12_V_0<A_SINT_CC_SCALbx24_waycap)) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0
              ]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) || (xpc10nz==10'd576/*US*/) || (xpc10nz==6'd37/*US*/)) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]==2'd2/*MS*/) || (((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==1'd1/*MS*/)? (xpc10nz==10'd565/*US*/): (xpc10nz
              ==10'd558/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/)) || (xpc10nz==10'd565/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [2'd2]!=0/*MS*/) || (xpc10nz==10'd540/*US*/) || (xpc10nz==6'd59/*US*/) || (xpc10nz==10'd571/*US*/) || ((xpc10nz==10'd558
              /*US*/) || (xpc10nz==10'd550/*US*/) || (xpc10nz==10'd565/*US*/)) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==2'd3/*MS*/)) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==2'd2/*MS*/);

               A_SINT_CC_MAPR10NoCE3_ARA0_WEN0 = ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==2'd3/*MS*/)? (((((xpc10nz==5'd20/*US*/) || (xpc10nz
              ==7'd65/*US*/) && (TCCl0_12_V_0<A_SINT_CC_SCALbx24_waycap)) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [0]!=2'd3/*MS*/) || (xpc10nz==6'd37/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/)) && (A_sA_SINT_CC_SCALbx20_ARA0
              [1'd1]!=2'd3/*MS*/) || (xpc10nz==10'd576/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) || (xpc10nz==10'd588/*US*/)) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) || (xpc10nz==10'd599/*US*/)) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) || 
              (xpc10nz==10'd609/*US*/) || (xpc10nz==6'd50/*US*/) || ((xpc10nz==10'd550/*US*/) || (xpc10nz==10'd558/*US*/) || (xpc10nz
              ==10'd565/*US*/)) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==2'd3/*MS*/): ((((((xpc10nz==5'd20/*US*/) || (xpc10nz==7'd65/*US*/) && 
              (TCCl0_12_V_0<A_SINT_CC_SCALbx24_waycap)) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]
              !=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [0]!=2'd3/*MS*/) || (xpc10nz==6'd37/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/)) && (A_sA_SINT_CC_SCALbx20_ARA0
              [1'd1]!=2'd3/*MS*/) || (xpc10nz==10'd576/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) || (xpc10nz==10'd588/*US*/)) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) || (xpc10nz==10'd599/*US*/)) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [1'd1]!=0/*MS*/) || ((xpc10nz==10'd609/*US*/) || (xpc10nz==6'd50/*US*/)) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/)) && (A_sA_SINT_CC_SCALbx20_ARA0
              [2'd3]==2'd3/*MS*/)) || ((TCin1_9_V_4==3'd4/*US*/)? !A_SINT_CC_MAPR10NoCE3_ARA0_RDD0 && (xpc10nz==9'd473/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [TCin1_9_V_4]==2'd3/*MS*/): ((((A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd3/*MS*/)? (xpc10nz==9'd503/*US*/) || (xpc10nz
              ==9'd259/*US*/): ((xpc10nz==9'd503/*US*/) || (xpc10nz==9'd259/*US*/)) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=0/*MS*/) && 
              (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd2/*MS*/)) || ((xpc10nz
              ==9'd503/*US*/) || (xpc10nz==9'd259/*US*/)) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==0/*MS*/) || ((xpc10nz==9'd503/*US*/) || 
              (xpc10nz==9'd259/*US*/)) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==1'd1/*MS*/) || ((xpc10nz==9'd503/*US*/) || (xpc10nz
              ==9'd259/*US*/)) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd2/*MS*/)) && (TCin1_9_V_4>=3'd4) || ((A_sA_SINT_CC_SCALbx22_ARB0
              [TCin1_9_V_4]==2'd3/*MS*/)? !A_SINT_CC_MAPR10NoCE3_ARA0_RDD0 && (xpc10nz==9'd473/*US*/): !A_SINT_CC_MAPR10NoCE3_ARA0_RDD0
               && (xpc10nz==9'd473/*US*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4
              ]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd2/*MS*/)) || !A_SINT_CC_MAPR10NoCE3_ARA0_RDD0 && (xpc10nz
              ==9'd473/*US*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==0/*MS*/) || !A_SINT_CC_MAPR10NoCE3_ARA0_RDD0 && (xpc10nz==
              9'd473/*US*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==1'd1/*MS*/) || !A_SINT_CC_MAPR10NoCE3_ARA0_RDD0 && (xpc10nz==
              9'd473/*US*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd2/*MS*/)) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd3
              /*MS*/)) || (TCCl0_12_V_1<3'd4) && (A_sA_SINT_CC_SCALbx20_ARA0[TCCl0_12_V_1]==2'd3/*MS*/) && (xpc10nz==10'd532/*US*/) || 
              (((A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]==2'd3/*MS*/)? 1'd1: (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim
              ]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim
              ]!=2'd2/*MS*/)) || (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]==0/*MS*/) || (A_sA_SINT_CC_SCALbx22_ARB0
              [A_SINT_CC_SCALbx24_next_victim]==1'd1/*MS*/) || (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]==2'd2/*MS*/)) && 
              (xpc10nz==9'd289/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]==2'd3/*MS*/) || ((xpc10nz==5'd20
              /*US*/) || (xpc10nz==7'd65/*US*/) && (TCCl0_12_V_0<A_SINT_CC_SCALbx24_waycap)) && (A_sA_SINT_CC_SCALbx20_ARA0[0]==2'd3/*MS*/) || 
              (((xpc10nz==5'd20/*US*/) || (xpc10nz==7'd65/*US*/) && (TCCl0_12_V_0<A_SINT_CC_SCALbx24_waycap)) && (A_sA_SINT_CC_SCALbx20_ARA0
              [0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [0]!=2'd3/*MS*/) || (xpc10nz==6'd37/*US*/)) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]==2'd3/*MS*/) || (((A_sA_SINT_CC_SCALbx20_ARA0
              [2'd2]==2'd2/*MS*/)? (xpc10nz==10'd558/*US*/) || (xpc10nz==10'd565/*US*/): (xpc10nz==10'd550/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/)) || ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==1'd1/*MS*/)? (xpc10nz
              ==10'd565/*US*/): (xpc10nz==10'd558/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/)) || (xpc10nz==10'd565/*US*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) || (xpc10nz==6'd59/*US*/) || (xpc10nz==10'd571/*US*/)) && (A_sA_SINT_CC_SCALbx20_ARA0
              [2'd3]==2'd3/*MS*/);

               end 
              
      case (xpc10nz) // synthesis full_case 
          5'd20/*US*/:  begin 
              if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==0/*MS*/) && !xpc10_stall
              )  begin 
                       A_SINT_CC_MAPR10NoCE0_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE0_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==1'd1/*MS*/) && 
              !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE1_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE1_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==2'd2/*MS*/) && 
              !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE2_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE2_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==2'd3/*MS*/) && 
              !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE3_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE3_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==0/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE0_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE0_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==1'd1/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE1_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE1_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==2'd2/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE2_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE2_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==2'd3/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE3_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE3_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]==0/*MS*/) && !xpc10_stall
              )  begin 
                       A_SINT_CC_MAPR10NoCE0_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE0_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]==1'd1/*MS*/) && !xpc10_stall
              )  begin 
                       A_SINT_CC_MAPR10NoCE1_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE1_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]==2'd2/*MS*/) && !xpc10_stall
              )  begin 
                       A_SINT_CC_MAPR10NoCE2_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE2_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]==2'd3/*MS*/) && !xpc10_stall
              )  begin 
                       A_SINT_CC_MAPR10NoCE3_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE3_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[0]==0/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE0_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE0_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[0]==1'd1/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE1_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE1_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[0]==2'd2/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE2_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE2_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[0]==2'd3/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE3_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE3_ARA0_AD0 = 13'd0;
                       end 
                       end 
              
          6'd37/*US*/:  begin 
              if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==0/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE0_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE0_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==1'd1/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE1_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE1_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==2'd2/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE2_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE2_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==2'd3/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE3_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE3_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==0/*MS*/) && !xpc10_stall
              )  begin 
                       A_SINT_CC_MAPR10NoCE0_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE0_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==1'd1/*MS*/) && 
              !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE1_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE1_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==2'd2/*MS*/) && 
              !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE2_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE2_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==2'd3/*MS*/) && 
              !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE3_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE3_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]==0/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE0_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE0_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]==1'd1/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE1_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE1_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]==2'd2/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE2_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE2_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]==2'd3/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE3_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE3_ARA0_AD0 = 13'd0;
                       end 
                       end 
              
          6'd50/*US*/:  begin 
              if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==0/*MS*/) && !xpc10_stall
              )  begin 
                       A_SINT_CC_MAPR10NoCE0_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE0_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==1'd1/*MS*/) && 
              !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE1_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE1_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==2'd2/*MS*/) && 
              !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE2_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE2_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==2'd3/*MS*/) && 
              !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE3_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE3_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==0/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE0_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE0_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==1'd1/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE1_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE1_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==2'd2/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE2_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE2_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==2'd3/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE3_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE3_ARA0_AD0 = 13'd0;
                       end 
                       end 
              endcase
      if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==0/*MS*/) && (xpc10nz==6'd59/*US*/) && !xpc10_stall)  begin 
               A_SINT_CC_MAPR10NoCE0_ARA0_WRD0 = 32'd0;
               A_SINT_CC_MAPR10NoCE0_ARA0_AD0 = 13'd0;
               end 
              if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==1'd1/*MS*/) && (xpc10nz==6'd59/*US*/) && !xpc10_stall)  begin 
               A_SINT_CC_MAPR10NoCE1_ARA0_WRD0 = 32'd0;
               A_SINT_CC_MAPR10NoCE1_ARA0_AD0 = 13'd0;
               end 
              
      case (xpc10nz) // synthesis full_case 
          6'd59/*US*/:  begin 
              if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==2'd2/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE2_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE2_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==2'd3/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE3_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE3_ARA0_AD0 = 13'd0;
                       end 
                       end 
              
          7'd65/*US*/:  begin 
              if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==0/*MS*/) && (TCCl0_12_V_0
              <A_SINT_CC_SCALbx24_waycap) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE0_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE0_ARA0_AD0 = TCCl0_12_V_0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==1'd1/*MS*/) && 
              (TCCl0_12_V_0<A_SINT_CC_SCALbx24_waycap) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE1_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE1_ARA0_AD0 = TCCl0_12_V_0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==2'd2/*MS*/) && 
              (TCCl0_12_V_0<A_SINT_CC_SCALbx24_waycap) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE2_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE2_ARA0_AD0 = TCCl0_12_V_0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==2'd3/*MS*/) && 
              (TCCl0_12_V_0<A_SINT_CC_SCALbx24_waycap) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE3_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE3_ARA0_AD0 = TCCl0_12_V_0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==0/*MS*/) && (TCCl0_12_V_0<A_SINT_CC_SCALbx24_waycap) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE0_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE0_ARA0_AD0 = TCCl0_12_V_0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==1'd1/*MS*/) && (TCCl0_12_V_0<A_SINT_CC_SCALbx24_waycap) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE1_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE1_ARA0_AD0 = TCCl0_12_V_0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==2'd2/*MS*/) && (TCCl0_12_V_0<A_SINT_CC_SCALbx24_waycap) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE2_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE2_ARA0_AD0 = TCCl0_12_V_0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==2'd3/*MS*/) && (TCCl0_12_V_0<A_SINT_CC_SCALbx24_waycap) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE3_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE3_ARA0_AD0 = TCCl0_12_V_0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]==0/*MS*/) && (TCCl0_12_V_0
              <A_SINT_CC_SCALbx24_waycap) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE0_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE0_ARA0_AD0 = TCCl0_12_V_0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]==1'd1/*MS*/) && (TCCl0_12_V_0
              <A_SINT_CC_SCALbx24_waycap) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE1_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE1_ARA0_AD0 = TCCl0_12_V_0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]==2'd2/*MS*/) && (TCCl0_12_V_0
              <A_SINT_CC_SCALbx24_waycap) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE2_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE2_ARA0_AD0 = TCCl0_12_V_0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]==2'd3/*MS*/) && (TCCl0_12_V_0
              <A_SINT_CC_SCALbx24_waycap) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE3_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE3_ARA0_AD0 = TCCl0_12_V_0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[0]==0/*MS*/) && (TCCl0_12_V_0<A_SINT_CC_SCALbx24_waycap) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE0_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE0_ARA0_AD0 = TCCl0_12_V_0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[0]==1'd1/*MS*/) && (TCCl0_12_V_0<A_SINT_CC_SCALbx24_waycap) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE1_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE1_ARA0_AD0 = TCCl0_12_V_0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[0]==2'd2/*MS*/) && (TCCl0_12_V_0<A_SINT_CC_SCALbx24_waycap) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE2_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE2_ARA0_AD0 = TCCl0_12_V_0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[0]==2'd3/*MS*/) && (TCCl0_12_V_0<A_SINT_CC_SCALbx24_waycap) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE3_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE3_ARA0_AD0 = TCCl0_12_V_0;
                       end 
                       end 
              endcase
      if ((TCha3_10_V_0>=0) && (xpc10nz==7'd106/*US*/) && !xpc10_stall)  begin 
               isMODULUS10_DD = A_SINT_CC_SCALbx24_waycap;
               isMODULUS10_NN = TCha3_10_V_0;
               end 
              if (!xpc10_stall) 
          case (xpc10nz) // synthesis full_case 
              8'd171/*US*/:  begin 
                   isMODULUS10_DD = A_SINT_CC_SCALbx24_waycap;
                   isMODULUS10_NN = TCha3_10_V_0;
                   end 
                  
              8'd236/*US*/:  begin 
                   A_SINT_CC_MAPR10NoCE3_ARA0_AD0 = TClo6_9_V_1;
                   A_SINT_CC_MAPR10NoCE2_ARA0_AD0 = TClo6_9_V_1;
                   A_SINT_CC_MAPR10NoCE1_ARA0_AD0 = TClo6_9_V_1;
                   A_SINT_CC_MAPR10NoCE0_ARA0_AD0 = TClo6_9_V_1;
                   end 
                  endcase
          if ((TClo6_9_V_0!=3'd4/*US*/) && (xpc10nz==8'd236/*US*/) && (TTMT4Main_V_11==((A_sA_SINT_CC_SCALbx20_ARA0[TClo6_9_V_0]==2'd3
      /*MS*/)? ((xpc10nz==8'd237/*US*/)? A_SINT_CC_MAPR10NoCE3_ARA0_RDD0: SINTCCMAPR10NoCE3ARA0RRh10hold): ((A_sA_SINT_CC_SCALbx20_ARA0
      [TClo6_9_V_0]==2'd2/*MS*/)? ((xpc10nz==8'd237/*US*/)? A_SINT_CC_MAPR10NoCE2_ARA0_RDD0: SINTCCMAPR10NoCE2ARA0RRh10hold): ((A_sA_SINT_CC_SCALbx20_ARA0
      [TClo6_9_V_0]==1'd1/*MS*/)? ((xpc10nz==8'd237/*US*/)? A_SINT_CC_MAPR10NoCE1_ARA0_RDD0: SINTCCMAPR10NoCE1ARA0RRh10hold): ((A_sA_SINT_CC_SCALbx20_ARA0
      [TClo6_9_V_0]==0/*MS*/)? ((xpc10nz==8'd237/*US*/)? A_SINT_CC_MAPR10NoCE0_ARA0_RDD0: SINTCCMAPR10NoCE0ARA0RRh10hold): 1'bx))))) && 
      !xpc10_stall)  begin 
               A_SINT_CC_MAPR12NoCE3_ARB0_AD0 = TClo6_9_V_1;
               A_SINT_CC_MAPR12NoCE2_ARB0_AD0 = TClo6_9_V_1;
               A_SINT_CC_MAPR12NoCE1_ARB0_AD0 = TClo6_9_V_1;
               A_SINT_CC_MAPR12NoCE0_ARB0_AD0 = TClo6_9_V_1;
               end 
              if (!xpc10_stall)  begin if ((xpc10nz==8'd239/*US*/))  A_64_US_CC_SCALbx26_ARA0_AD0 = TClo6_9_V_2;
               end 
          if ((TClo6_9_V_0>=3'd4) && (TClo6_9_V_0!=3'd4/*US*/) && (xpc10nz==8'd242/*US*/) && !xpc10_stall)  begin 
               A_SINT_CC_MAPR12NoCE3_ARB0_AD0 = TClo6_9_V_1;
               A_SINT_CC_MAPR12NoCE2_ARB0_AD0 = TClo6_9_V_1;
               A_SINT_CC_MAPR12NoCE1_ARB0_AD0 = TClo6_9_V_1;
               A_SINT_CC_MAPR12NoCE0_ARB0_AD0 = TClo6_9_V_1;
               end 
              if ((xpc10nz==8'd255/*US*/) && !xpc10_stall)  begin 
               A_64_US_CC_SCALbx26_ARA0_WRD0 = TTMT4Main_V_6;
               A_64_US_CC_SCALbx26_ARA0_AD0 = 32'hffffffff&TCin1_9_V_3;
               end 
              if ((xpc10nz==9'd259/*US*/))  begin 
              if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4
              ]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==0/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR12NoCE0_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE0_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd3/*MS*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [TCin1_9_V_4]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==1'd1/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR12NoCE1_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE1_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd3/*MS*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [TCin1_9_V_4]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd2/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR12NoCE2_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE2_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd3/*MS*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [TCin1_9_V_4]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd3/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR12NoCE3_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE3_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
              [TCin1_9_V_4]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4
              ]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=0/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE0_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE0_ARA0_AD0 = TCin1_9_V_5;
                       end 
                      if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
              [TCin1_9_V_4]==0/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE0_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE0_ARA0_AD0 = TCin1_9_V_5;
                       A_SINT_CC_MAPR12NoCE0_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE0_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
              [TCin1_9_V_4]==1'd1/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE0_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE0_ARA0_AD0 = TCin1_9_V_5;
                       A_SINT_CC_MAPR12NoCE1_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE1_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
              [TCin1_9_V_4]==2'd2/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE0_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE0_ARA0_AD0 = TCin1_9_V_5;
                       A_SINT_CC_MAPR12NoCE2_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE2_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
              [TCin1_9_V_4]==2'd3/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE0_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE0_ARA0_AD0 = TCin1_9_V_5;
                       A_SINT_CC_MAPR12NoCE3_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE3_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==1'd1/*MS*/) && 
              (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
              [TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=0/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE1_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE1_ARA0_AD0 = TCin1_9_V_5;
                       end 
                      if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==1'd1/*MS*/) && 
              (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==0/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE1_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE1_ARA0_AD0 = TCin1_9_V_5;
                       A_SINT_CC_MAPR12NoCE0_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE0_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==1'd1/*MS*/) && 
              (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==1'd1/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE1_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE1_ARA0_AD0 = TCin1_9_V_5;
                       A_SINT_CC_MAPR12NoCE1_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE1_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==1'd1/*MS*/) && 
              (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd2/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE1_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE1_ARA0_AD0 = TCin1_9_V_5;
                       A_SINT_CC_MAPR12NoCE2_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE2_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==1'd1/*MS*/) && 
              (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd3/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE1_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE1_ARA0_AD0 = TCin1_9_V_5;
                       A_SINT_CC_MAPR12NoCE3_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE3_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd2/*MS*/) && 
              (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
              [TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=0/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE2_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE2_ARA0_AD0 = TCin1_9_V_5;
                       end 
                      if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd2/*MS*/) && 
              (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==0/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE2_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE2_ARA0_AD0 = TCin1_9_V_5;
                       A_SINT_CC_MAPR12NoCE0_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE0_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd2/*MS*/) && 
              (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==1'd1/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE2_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE2_ARA0_AD0 = TCin1_9_V_5;
                       A_SINT_CC_MAPR12NoCE1_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE1_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd2/*MS*/) && 
              (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd2/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE2_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE2_ARA0_AD0 = TCin1_9_V_5;
                       A_SINT_CC_MAPR12NoCE2_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE2_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd2/*MS*/) && 
              (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd3/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE2_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE2_ARA0_AD0 = TCin1_9_V_5;
                       A_SINT_CC_MAPR12NoCE3_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE3_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd3/*MS*/) && 
              (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
              [TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=0/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE3_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE3_ARA0_AD0 = TCin1_9_V_5;
                       end 
                      if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd3/*MS*/) && 
              (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==0/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE3_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE3_ARA0_AD0 = TCin1_9_V_5;
                       A_SINT_CC_MAPR12NoCE0_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE0_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd3/*MS*/) && 
              (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==1'd1/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE3_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE3_ARA0_AD0 = TCin1_9_V_5;
                       A_SINT_CC_MAPR12NoCE1_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE1_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd3/*MS*/) && 
              (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd2/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE3_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE3_ARA0_AD0 = TCin1_9_V_5;
                       A_SINT_CC_MAPR12NoCE2_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE2_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd3/*MS*/) && 
              (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd3/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE3_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE3_ARA0_AD0 = TCin1_9_V_5;
                       A_SINT_CC_MAPR12NoCE3_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE3_ARB0_AD0 = TCin1_9_V_5;
                       end 
                       end 
              if (!xpc10_stall) 
          case (xpc10nz) // synthesis full_case 
              9'd285/*US*/:  begin 
                   A_SINT_CC_MAPR10NoCE3_ARA0_AD0 = TCin1_9_V_5;
                   A_SINT_CC_MAPR10NoCE2_ARA0_AD0 = TCin1_9_V_5;
                   A_SINT_CC_MAPR10NoCE1_ARA0_AD0 = TCin1_9_V_5;
                   A_SINT_CC_MAPR10NoCE0_ARA0_AD0 = TCin1_9_V_5;
                   end 
                  
              9'd287/*US*/:  begin 
                   A_SINT_CC_MAPR12NoCE3_ARB0_AD0 = TCin1_9_V_5;
                   A_SINT_CC_MAPR12NoCE2_ARB0_AD0 = TCin1_9_V_5;
                   A_SINT_CC_MAPR12NoCE1_ARB0_AD0 = TCin1_9_V_5;
                   A_SINT_CC_MAPR12NoCE0_ARB0_AD0 = TCin1_9_V_5;
                   end 
                  endcase
          if ((xpc10nz==9'd289/*US*/))  begin 
              if ((A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim
              ]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [A_SINT_CC_SCALbx24_next_victim]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]==0/*MS*/) && 
              !xpc10_stall)  begin 
                       A_SINT_CC_MAPR12NoCE0_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE0_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim
              ]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [A_SINT_CC_SCALbx24_next_victim]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]==1'd1/*MS*/) && 
              !xpc10_stall)  begin 
                       A_SINT_CC_MAPR12NoCE1_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE1_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim
              ]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [A_SINT_CC_SCALbx24_next_victim]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]==2'd2/*MS*/) && 
              !xpc10_stall)  begin 
                       A_SINT_CC_MAPR12NoCE2_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE2_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim
              ]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [A_SINT_CC_SCALbx24_next_victim]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]==2'd3/*MS*/) && 
              !xpc10_stall)  begin 
                       A_SINT_CC_MAPR12NoCE3_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE3_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]==0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim
              ]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
              [A_SINT_CC_SCALbx24_next_victim]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]!=0/*MS*/) && 
              !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE0_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE0_ARA0_AD0 = TCin1_9_V_5;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]==0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim
              ]==0/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE0_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE0_ARA0_AD0 = TCin1_9_V_5;
                       A_SINT_CC_MAPR12NoCE0_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE0_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]==0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim
              ]==1'd1/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE0_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE0_ARA0_AD0 = TCin1_9_V_5;
                       A_SINT_CC_MAPR12NoCE1_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE1_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]==0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim
              ]==2'd2/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE0_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE0_ARA0_AD0 = TCin1_9_V_5;
                       A_SINT_CC_MAPR12NoCE2_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE2_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]==0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim
              ]==2'd3/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE0_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE0_ARA0_AD0 = TCin1_9_V_5;
                       A_SINT_CC_MAPR12NoCE3_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE3_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]==1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim
              ]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
              [A_SINT_CC_SCALbx24_next_victim]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]!=0/*MS*/) && 
              !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE1_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE1_ARA0_AD0 = TCin1_9_V_5;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]==1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim
              ]==0/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE1_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE1_ARA0_AD0 = TCin1_9_V_5;
                       A_SINT_CC_MAPR12NoCE0_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE0_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]==1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim
              ]==1'd1/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE1_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE1_ARA0_AD0 = TCin1_9_V_5;
                       A_SINT_CC_MAPR12NoCE1_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE1_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]==1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim
              ]==2'd2/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE1_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE1_ARA0_AD0 = TCin1_9_V_5;
                       A_SINT_CC_MAPR12NoCE2_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE2_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]==1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim
              ]==2'd3/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE1_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE1_ARA0_AD0 = TCin1_9_V_5;
                       A_SINT_CC_MAPR12NoCE3_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE3_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]==2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim
              ]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
              [A_SINT_CC_SCALbx24_next_victim]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]!=0/*MS*/) && 
              !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE2_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE2_ARA0_AD0 = TCin1_9_V_5;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]==2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim
              ]==0/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE2_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE2_ARA0_AD0 = TCin1_9_V_5;
                       A_SINT_CC_MAPR12NoCE0_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE0_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]==2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim
              ]==1'd1/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE2_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE2_ARA0_AD0 = TCin1_9_V_5;
                       A_SINT_CC_MAPR12NoCE1_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE1_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]==2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim
              ]==2'd2/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE2_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE2_ARA0_AD0 = TCin1_9_V_5;
                       A_SINT_CC_MAPR12NoCE2_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE2_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]==2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim
              ]==2'd3/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE2_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE2_ARA0_AD0 = TCin1_9_V_5;
                       A_SINT_CC_MAPR12NoCE3_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE3_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]==2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim
              ]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
              [A_SINT_CC_SCALbx24_next_victim]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]!=0/*MS*/) && 
              !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE3_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE3_ARA0_AD0 = TCin1_9_V_5;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]==2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim
              ]==0/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE3_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE3_ARA0_AD0 = TCin1_9_V_5;
                       A_SINT_CC_MAPR12NoCE0_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE0_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]==2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim
              ]==1'd1/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE3_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE3_ARA0_AD0 = TCin1_9_V_5;
                       A_SINT_CC_MAPR12NoCE1_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE1_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]==2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim
              ]==2'd2/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE3_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE3_ARA0_AD0 = TCin1_9_V_5;
                       A_SINT_CC_MAPR12NoCE2_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE2_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]==2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim
              ]==2'd3/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE3_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE3_ARA0_AD0 = TCin1_9_V_5;
                       A_SINT_CC_MAPR12NoCE3_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE3_ARB0_AD0 = TCin1_9_V_5;
                       end 
                       end 
              if ((A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]==0/*MS*/) && (xpc10nz==9'd314/*US*/) && !xpc10_stall)  begin 
               A_SINT_CC_MAPR12NoCE0_ARB0_WRD0 = TCin1_9_V_2;
               A_SINT_CC_MAPR12NoCE0_ARB0_AD0 = TCin1_9_V_5;
               end 
              if ((xpc10nz==9'd314/*US*/))  begin 
              if ((A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]==1'd1/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR12NoCE1_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE1_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if ((A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]==2'd2/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR12NoCE2_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE2_ARB0_AD0 = TCin1_9_V_5;
                       end 
                       end 
              if ((A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]==0/*MS*/) && (xpc10nz==9'd324/*US*/) && !xpc10_stall)  begin 
               A_SINT_CC_MAPR12NoCE0_ARB0_WRD0 = TCin1_9_V_2;
               A_SINT_CC_MAPR12NoCE0_ARB0_AD0 = TCin1_9_V_5;
               end 
              if ((A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]==1'd1/*MS*/) && (xpc10nz==9'd324/*US*/) && !xpc10_stall
      )  begin 
               A_SINT_CC_MAPR12NoCE1_ARB0_WRD0 = TCin1_9_V_2;
               A_SINT_CC_MAPR12NoCE1_ARB0_AD0 = TCin1_9_V_5;
               end 
              if ((A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]==0/*MS*/) && (xpc10nz==9'd327/*US*/) && !xpc10_stall)  begin 
               A_SINT_CC_MAPR12NoCE0_ARB0_WRD0 = TCin1_9_V_2;
               A_SINT_CC_MAPR12NoCE0_ARB0_AD0 = TCin1_9_V_5;
               end 
              if ((A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==0/*MS*/) && (xpc10nz==9'd330/*US*/) && !xpc10_stall)  begin 
               A_SINT_CC_MAPR12NoCE0_ARB0_WRD0 = TCin1_9_V_2;
               A_SINT_CC_MAPR12NoCE0_ARB0_AD0 = TCin1_9_V_5;
               end 
              if ((xpc10nz==9'd330/*US*/))  begin 
              if ((A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==1'd1/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR12NoCE1_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE1_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if ((A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd2/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR12NoCE2_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE2_ARB0_AD0 = TCin1_9_V_5;
                       end 
                       end 
              if ((A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==0/*MS*/) && (xpc10nz==9'd335/*US*/) && !xpc10_stall)  begin 
               A_SINT_CC_MAPR12NoCE0_ARB0_WRD0 = TCin1_9_V_2;
               A_SINT_CC_MAPR12NoCE0_ARB0_AD0 = TCin1_9_V_5;
               end 
              if ((A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==1'd1/*MS*/) && (xpc10nz==9'd335/*US*/) && !xpc10_stall)  begin 
               A_SINT_CC_MAPR12NoCE1_ARB0_WRD0 = TCin1_9_V_2;
               A_SINT_CC_MAPR12NoCE1_ARB0_AD0 = TCin1_9_V_5;
               end 
              if ((A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==0/*MS*/) && (xpc10nz==9'd338/*US*/) && !xpc10_stall)  begin 
               A_SINT_CC_MAPR12NoCE0_ARB0_WRD0 = TCin1_9_V_2;
               A_SINT_CC_MAPR12NoCE0_ARB0_AD0 = TCin1_9_V_5;
               end 
              if ((TCha6_10_V_0>=0) && (xpc10nz==9'd342/*US*/) && !xpc10_stall)  begin 
               isMODULUS10_DD = A_SINT_CC_SCALbx24_waycap;
               isMODULUS10_NN = TCha6_10_V_0;
               end 
              if (!xpc10_stall) 
          case (xpc10nz) // synthesis full_case 
              9'd407/*US*/:  begin 
                   isMODULUS10_DD = A_SINT_CC_SCALbx24_waycap;
                   isMODULUS10_NN = TCha6_10_V_0;
                   end 
                  
              9'd472/*US*/:  begin 
                   A_SINT_CC_MAPR10NoCE3_ARA0_AD0 = TCin1_9_V_5;
                   A_SINT_CC_MAPR10NoCE2_ARA0_AD0 = TCin1_9_V_5;
                   A_SINT_CC_MAPR10NoCE1_ARA0_AD0 = TCin1_9_V_5;
                   A_SINT_CC_MAPR10NoCE0_ARA0_AD0 = TCin1_9_V_5;
                   end 
                  endcase
          
      case (xpc10nz) // synthesis full_case 
          9'd473/*US*/:  begin 
              if ((TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4
              ]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=0/*MS*/) && 
              (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==0/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR12NoCE0_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE0_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if ((TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4
              ]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==1'd1/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR12NoCE1_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE1_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if ((TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4
              ]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd2/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR12NoCE2_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE2_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if ((TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4
              ]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd3/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR12NoCE3_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE3_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if (((xpc10nz==9'd473/*US*/)? !A_SINT_CC_MAPR10NoCE0_ARA0_RDD0 && !xpc10_stall: !SINTCCMAPR10NoCE0ARA0RRh10hold
               && !xpc10_stall) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=1'd1
              /*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd3/*MS*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==0/*MS*/) && (TCin1_9_V_4!=3'd4/*US*/))  begin 
                       A_SINT_CC_MAPR10NoCE0_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE0_ARA0_AD0 = TCin1_9_V_5;
                       end 
                      if (((xpc10nz==9'd473/*US*/)? !A_SINT_CC_MAPR10NoCE0_ARA0_RDD0 && !xpc10_stall: !SINTCCMAPR10NoCE0ARA0RRh10hold
               && !xpc10_stall) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==0/*MS*/) && 
              (TCin1_9_V_4!=3'd4/*US*/))  begin 
                       A_SINT_CC_MAPR10NoCE0_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE0_ARA0_AD0 = TCin1_9_V_5;
                       A_SINT_CC_MAPR12NoCE0_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE0_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if (((xpc10nz==9'd473/*US*/)? !A_SINT_CC_MAPR10NoCE0_ARA0_RDD0 && !xpc10_stall: !SINTCCMAPR10NoCE0ARA0RRh10hold
               && !xpc10_stall) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==
              0/*MS*/) && (TCin1_9_V_4!=3'd4/*US*/))  begin 
                       A_SINT_CC_MAPR10NoCE0_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE0_ARA0_AD0 = TCin1_9_V_5;
                       A_SINT_CC_MAPR12NoCE1_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE1_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if (((xpc10nz==9'd473/*US*/)? !A_SINT_CC_MAPR10NoCE0_ARA0_RDD0 && !xpc10_stall: !SINTCCMAPR10NoCE0ARA0RRh10hold
               && !xpc10_stall) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==
              0/*MS*/) && (TCin1_9_V_4!=3'd4/*US*/))  begin 
                       A_SINT_CC_MAPR10NoCE0_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE0_ARA0_AD0 = TCin1_9_V_5;
                       A_SINT_CC_MAPR12NoCE2_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE2_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if (((xpc10nz==9'd473/*US*/)? !A_SINT_CC_MAPR10NoCE0_ARA0_RDD0 && !xpc10_stall: !SINTCCMAPR10NoCE0ARA0RRh10hold
               && !xpc10_stall) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==
              0/*MS*/) && (TCin1_9_V_4!=3'd4/*US*/))  begin 
                       A_SINT_CC_MAPR10NoCE0_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE0_ARA0_AD0 = TCin1_9_V_5;
                       A_SINT_CC_MAPR12NoCE3_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE3_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if (((xpc10nz==9'd473/*US*/)? !A_SINT_CC_MAPR10NoCE0_ARA0_RDD0 && !xpc10_stall: !SINTCCMAPR10NoCE0ARA0RRh10hold
               && !xpc10_stall) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==0/*MS*/) && (TCin1_9_V_4==3'd4/*US*/))  begin 
                       A_SINT_CC_MAPR10NoCE0_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE0_ARA0_AD0 = TCin1_9_V_5;
                       end 
                      if (((xpc10nz==9'd473/*US*/)? !A_SINT_CC_MAPR10NoCE1_ARA0_RDD0 && !xpc10_stall: !SINTCCMAPR10NoCE1ARA0RRh10hold
               && !xpc10_stall) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=1'd1
              /*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd3/*MS*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==1'd1/*MS*/) && (TCin1_9_V_4!=3'd4/*US*/))  begin 
                       A_SINT_CC_MAPR10NoCE1_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE1_ARA0_AD0 = TCin1_9_V_5;
                       end 
                      if (((xpc10nz==9'd473/*US*/)? !A_SINT_CC_MAPR10NoCE1_ARA0_RDD0 && !xpc10_stall: !SINTCCMAPR10NoCE1ARA0RRh10hold
               && !xpc10_stall) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==1'd1
              /*MS*/) && (TCin1_9_V_4!=3'd4/*US*/))  begin 
                       A_SINT_CC_MAPR10NoCE1_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE1_ARA0_AD0 = TCin1_9_V_5;
                       A_SINT_CC_MAPR12NoCE0_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE0_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if (((xpc10nz==9'd473/*US*/)? !A_SINT_CC_MAPR10NoCE1_ARA0_RDD0 && !xpc10_stall: !SINTCCMAPR10NoCE1ARA0RRh10hold
               && !xpc10_stall) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==
              1'd1/*MS*/) && (TCin1_9_V_4!=3'd4/*US*/))  begin 
                       A_SINT_CC_MAPR10NoCE1_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE1_ARA0_AD0 = TCin1_9_V_5;
                       A_SINT_CC_MAPR12NoCE1_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE1_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if (((xpc10nz==9'd473/*US*/)? !A_SINT_CC_MAPR10NoCE1_ARA0_RDD0 && !xpc10_stall: !SINTCCMAPR10NoCE1ARA0RRh10hold
               && !xpc10_stall) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==
              1'd1/*MS*/) && (TCin1_9_V_4!=3'd4/*US*/))  begin 
                       A_SINT_CC_MAPR10NoCE1_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE1_ARA0_AD0 = TCin1_9_V_5;
                       A_SINT_CC_MAPR12NoCE2_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE2_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if (((xpc10nz==9'd473/*US*/)? !A_SINT_CC_MAPR10NoCE1_ARA0_RDD0 && !xpc10_stall: !SINTCCMAPR10NoCE1ARA0RRh10hold
               && !xpc10_stall) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==
              1'd1/*MS*/) && (TCin1_9_V_4!=3'd4/*US*/))  begin 
                       A_SINT_CC_MAPR10NoCE1_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE1_ARA0_AD0 = TCin1_9_V_5;
                       A_SINT_CC_MAPR12NoCE3_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE3_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if (((xpc10nz==9'd473/*US*/)? !A_SINT_CC_MAPR10NoCE1_ARA0_RDD0 && !xpc10_stall: !SINTCCMAPR10NoCE1ARA0RRh10hold
               && !xpc10_stall) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==1'd1/*MS*/) && (TCin1_9_V_4==3'd4/*US*/))  begin 
                       A_SINT_CC_MAPR10NoCE1_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE1_ARA0_AD0 = TCin1_9_V_5;
                       end 
                      if (((xpc10nz==9'd473/*US*/)? !A_SINT_CC_MAPR10NoCE2_ARA0_RDD0 && !xpc10_stall: !SINTCCMAPR10NoCE2ARA0RRh10hold
               && !xpc10_stall) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=1'd1
              /*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd3/*MS*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd2/*MS*/) && (TCin1_9_V_4!=3'd4/*US*/))  begin 
                       A_SINT_CC_MAPR10NoCE2_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE2_ARA0_AD0 = TCin1_9_V_5;
                       end 
                      if (((xpc10nz==9'd473/*US*/)? !A_SINT_CC_MAPR10NoCE2_ARA0_RDD0 && !xpc10_stall: !SINTCCMAPR10NoCE2ARA0RRh10hold
               && !xpc10_stall) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd2
              /*MS*/) && (TCin1_9_V_4!=3'd4/*US*/))  begin 
                       A_SINT_CC_MAPR10NoCE2_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE2_ARA0_AD0 = TCin1_9_V_5;
                       A_SINT_CC_MAPR12NoCE0_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE0_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if (((xpc10nz==9'd473/*US*/)? !A_SINT_CC_MAPR10NoCE2_ARA0_RDD0 && !xpc10_stall: !SINTCCMAPR10NoCE2ARA0RRh10hold
               && !xpc10_stall) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==
              2'd2/*MS*/) && (TCin1_9_V_4!=3'd4/*US*/))  begin 
                       A_SINT_CC_MAPR10NoCE2_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE2_ARA0_AD0 = TCin1_9_V_5;
                       A_SINT_CC_MAPR12NoCE1_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE1_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if (((xpc10nz==9'd473/*US*/)? !A_SINT_CC_MAPR10NoCE2_ARA0_RDD0 && !xpc10_stall: !SINTCCMAPR10NoCE2ARA0RRh10hold
               && !xpc10_stall) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==
              2'd2/*MS*/) && (TCin1_9_V_4!=3'd4/*US*/))  begin 
                       A_SINT_CC_MAPR10NoCE2_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE2_ARA0_AD0 = TCin1_9_V_5;
                       A_SINT_CC_MAPR12NoCE2_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE2_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if (((xpc10nz==9'd473/*US*/)? !A_SINT_CC_MAPR10NoCE2_ARA0_RDD0 && !xpc10_stall: !SINTCCMAPR10NoCE2ARA0RRh10hold
               && !xpc10_stall) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==
              2'd2/*MS*/) && (TCin1_9_V_4!=3'd4/*US*/))  begin 
                       A_SINT_CC_MAPR10NoCE2_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE2_ARA0_AD0 = TCin1_9_V_5;
                       A_SINT_CC_MAPR12NoCE3_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE3_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if (((xpc10nz==9'd473/*US*/)? !A_SINT_CC_MAPR10NoCE2_ARA0_RDD0 && !xpc10_stall: !SINTCCMAPR10NoCE2ARA0RRh10hold
               && !xpc10_stall) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd2/*MS*/) && (TCin1_9_V_4==3'd4/*US*/))  begin 
                       A_SINT_CC_MAPR10NoCE2_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE2_ARA0_AD0 = TCin1_9_V_5;
                       end 
                      if (((xpc10nz==9'd473/*US*/)? !A_SINT_CC_MAPR10NoCE3_ARA0_RDD0 && !xpc10_stall: !SINTCCMAPR10NoCE3ARA0RRh10hold
               && !xpc10_stall) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=1'd1
              /*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd3/*MS*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd3/*MS*/) && (TCin1_9_V_4!=3'd4/*US*/))  begin 
                       A_SINT_CC_MAPR10NoCE3_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE3_ARA0_AD0 = TCin1_9_V_5;
                       end 
                      if (((xpc10nz==9'd473/*US*/)? !A_SINT_CC_MAPR10NoCE3_ARA0_RDD0 && !xpc10_stall: !SINTCCMAPR10NoCE3ARA0RRh10hold
               && !xpc10_stall) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd3
              /*MS*/) && (TCin1_9_V_4!=3'd4/*US*/))  begin 
                       A_SINT_CC_MAPR10NoCE3_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE3_ARA0_AD0 = TCin1_9_V_5;
                       A_SINT_CC_MAPR12NoCE0_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE0_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if (((xpc10nz==9'd473/*US*/)? !A_SINT_CC_MAPR10NoCE3_ARA0_RDD0 && !xpc10_stall: !SINTCCMAPR10NoCE3ARA0RRh10hold
               && !xpc10_stall) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==
              2'd3/*MS*/) && (TCin1_9_V_4!=3'd4/*US*/))  begin 
                       A_SINT_CC_MAPR10NoCE3_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE3_ARA0_AD0 = TCin1_9_V_5;
                       A_SINT_CC_MAPR12NoCE1_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE1_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if (((xpc10nz==9'd473/*US*/)? !A_SINT_CC_MAPR10NoCE3_ARA0_RDD0 && !xpc10_stall: !SINTCCMAPR10NoCE3ARA0RRh10hold
               && !xpc10_stall) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==
              2'd3/*MS*/) && (TCin1_9_V_4!=3'd4/*US*/))  begin 
                       A_SINT_CC_MAPR10NoCE3_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE3_ARA0_AD0 = TCin1_9_V_5;
                       A_SINT_CC_MAPR12NoCE2_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE2_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if (((xpc10nz==9'd473/*US*/)? !A_SINT_CC_MAPR10NoCE3_ARA0_RDD0 && !xpc10_stall: !SINTCCMAPR10NoCE3ARA0RRh10hold
               && !xpc10_stall) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==
              2'd3/*MS*/) && (TCin1_9_V_4!=3'd4/*US*/))  begin 
                       A_SINT_CC_MAPR10NoCE3_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE3_ARA0_AD0 = TCin1_9_V_5;
                       A_SINT_CC_MAPR12NoCE3_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE3_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if (((xpc10nz==9'd473/*US*/)? !A_SINT_CC_MAPR10NoCE3_ARA0_RDD0 && !xpc10_stall: !SINTCCMAPR10NoCE3ARA0RRh10hold
               && !xpc10_stall) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd3/*MS*/) && (TCin1_9_V_4==3'd4/*US*/))  begin 
                       A_SINT_CC_MAPR10NoCE3_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE3_ARA0_AD0 = TCin1_9_V_5;
                       end 
                       end 
              
          9'd503/*US*/:  begin 
              if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4
              ]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==0/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR12NoCE0_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE0_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd3/*MS*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [TCin1_9_V_4]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==1'd1/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR12NoCE1_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE1_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd3/*MS*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [TCin1_9_V_4]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd2/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR12NoCE2_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE2_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd3/*MS*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [TCin1_9_V_4]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd3/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR12NoCE3_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE3_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
              [TCin1_9_V_4]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4
              ]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=0/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE0_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE0_ARA0_AD0 = TCin1_9_V_5;
                       end 
                      if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
              [TCin1_9_V_4]==0/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE0_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE0_ARA0_AD0 = TCin1_9_V_5;
                       A_SINT_CC_MAPR12NoCE0_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE0_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
              [TCin1_9_V_4]==1'd1/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE0_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE0_ARA0_AD0 = TCin1_9_V_5;
                       A_SINT_CC_MAPR12NoCE1_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE1_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
              [TCin1_9_V_4]==2'd2/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE0_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE0_ARA0_AD0 = TCin1_9_V_5;
                       A_SINT_CC_MAPR12NoCE2_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE2_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
              [TCin1_9_V_4]==2'd3/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE0_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE0_ARA0_AD0 = TCin1_9_V_5;
                       A_SINT_CC_MAPR12NoCE3_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE3_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==1'd1/*MS*/) && 
              (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
              [TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=0/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE1_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE1_ARA0_AD0 = TCin1_9_V_5;
                       end 
                      if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==1'd1/*MS*/) && 
              (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==0/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE1_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE1_ARA0_AD0 = TCin1_9_V_5;
                       A_SINT_CC_MAPR12NoCE0_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE0_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==1'd1/*MS*/) && 
              (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==1'd1/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE1_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE1_ARA0_AD0 = TCin1_9_V_5;
                       A_SINT_CC_MAPR12NoCE1_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE1_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==1'd1/*MS*/) && 
              (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd2/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE1_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE1_ARA0_AD0 = TCin1_9_V_5;
                       A_SINT_CC_MAPR12NoCE2_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE2_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==1'd1/*MS*/) && 
              (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd3/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE1_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE1_ARA0_AD0 = TCin1_9_V_5;
                       A_SINT_CC_MAPR12NoCE3_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE3_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd2/*MS*/) && 
              (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
              [TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=0/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE2_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE2_ARA0_AD0 = TCin1_9_V_5;
                       end 
                      if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd2/*MS*/) && 
              (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==0/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE2_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE2_ARA0_AD0 = TCin1_9_V_5;
                       A_SINT_CC_MAPR12NoCE0_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE0_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd2/*MS*/) && 
              (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==1'd1/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE2_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE2_ARA0_AD0 = TCin1_9_V_5;
                       A_SINT_CC_MAPR12NoCE1_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE1_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd2/*MS*/) && 
              (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd2/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE2_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE2_ARA0_AD0 = TCin1_9_V_5;
                       A_SINT_CC_MAPR12NoCE2_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE2_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd2/*MS*/) && 
              (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd3/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE2_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE2_ARA0_AD0 = TCin1_9_V_5;
                       A_SINT_CC_MAPR12NoCE3_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE3_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd3/*MS*/) && 
              (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
              [TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=0/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE3_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE3_ARA0_AD0 = TCin1_9_V_5;
                       end 
                      if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd3/*MS*/) && 
              (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==0/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE3_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE3_ARA0_AD0 = TCin1_9_V_5;
                       A_SINT_CC_MAPR12NoCE0_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE0_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd3/*MS*/) && 
              (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==1'd1/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE3_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE3_ARA0_AD0 = TCin1_9_V_5;
                       A_SINT_CC_MAPR12NoCE1_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE1_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd3/*MS*/) && 
              (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd2/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE3_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE3_ARA0_AD0 = TCin1_9_V_5;
                       A_SINT_CC_MAPR12NoCE2_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE2_ARB0_AD0 = TCin1_9_V_5;
                       end 
                      if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd3/*MS*/) && 
              (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd3/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE3_ARA0_WRD0 = TCin1_9_V_0;
                       A_SINT_CC_MAPR10NoCE3_ARA0_AD0 = TCin1_9_V_5;
                       A_SINT_CC_MAPR12NoCE3_ARB0_WRD0 = TCin1_9_V_2;
                       A_SINT_CC_MAPR12NoCE3_ARB0_AD0 = TCin1_9_V_5;
                       end 
                       end 
              endcase
      if ((A_sA_SINT_CC_SCALbx20_ARA0[TCCl0_12_V_1]==0/*MS*/) && (xpc10nz==10'd528/*US*/) && !xpc10_stall)  begin 
               A_SINT_CC_MAPR10NoCE0_ARA0_WRD0 = 32'd0;
               A_SINT_CC_MAPR10NoCE0_ARA0_AD0 = TCCl0_12_V_0;
               end 
              
      case (xpc10nz) // synthesis full_case 
          10'd528/*US*/:  begin 
              if ((A_sA_SINT_CC_SCALbx20_ARA0[TCCl0_12_V_1]==1'd1/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE1_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE1_ARA0_AD0 = TCCl0_12_V_0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[TCCl0_12_V_1]==2'd2/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE2_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE2_ARA0_AD0 = TCCl0_12_V_0;
                       end 
                       end 
              
          10'd532/*US*/:  begin 
              if ((TCCl0_12_V_1<3'd4) && (A_sA_SINT_CC_SCALbx20_ARA0[TCCl0_12_V_1]==2'd3/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE3_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE3_ARA0_AD0 = TCCl0_12_V_0;
                       end 
                      if ((TCCl0_12_V_1<3'd4) && (A_sA_SINT_CC_SCALbx20_ARA0[TCCl0_12_V_1]==2'd2/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE2_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE2_ARA0_AD0 = TCCl0_12_V_0;
                       end 
                      if ((TCCl0_12_V_1<3'd4) && (A_sA_SINT_CC_SCALbx20_ARA0[TCCl0_12_V_1]==1'd1/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE1_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE1_ARA0_AD0 = TCCl0_12_V_0;
                       end 
                      if ((TCCl0_12_V_1<3'd4) && (A_sA_SINT_CC_SCALbx20_ARA0[TCCl0_12_V_1]==0/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE0_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE0_ARA0_AD0 = TCCl0_12_V_0;
                       end 
                       end 
              endcase
      if ((A_sA_SINT_CC_SCALbx20_ARA0[TCCl0_12_V_1]==0/*MS*/) && (xpc10nz==10'd534/*US*/) && !xpc10_stall)  begin 
               A_SINT_CC_MAPR10NoCE0_ARA0_WRD0 = 32'd0;
               A_SINT_CC_MAPR10NoCE0_ARA0_AD0 = TCCl0_12_V_0;
               end 
              if ((A_sA_SINT_CC_SCALbx20_ARA0[TCCl0_12_V_1]==1'd1/*MS*/) && (xpc10nz==10'd534/*US*/) && !xpc10_stall)  begin 
               A_SINT_CC_MAPR10NoCE1_ARA0_WRD0 = 32'd0;
               A_SINT_CC_MAPR10NoCE1_ARA0_AD0 = TCCl0_12_V_0;
               end 
              if ((A_sA_SINT_CC_SCALbx20_ARA0[TCCl0_12_V_1]==0/*MS*/) && (xpc10nz==10'd537/*US*/) && !xpc10_stall)  begin 
               A_SINT_CC_MAPR10NoCE0_ARA0_WRD0 = 32'd0;
               A_SINT_CC_MAPR10NoCE0_ARA0_AD0 = TCCl0_12_V_0;
               end 
              if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==0/*MS*/) && (xpc10nz==10'd540/*US*/) && !xpc10_stall)  begin 
               A_SINT_CC_MAPR10NoCE0_ARA0_WRD0 = 32'd0;
               A_SINT_CC_MAPR10NoCE0_ARA0_AD0 = 13'd0;
               end 
              if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==1'd1/*MS*/) && (xpc10nz==10'd540/*US*/) && !xpc10_stall)  begin 
               A_SINT_CC_MAPR10NoCE1_ARA0_WRD0 = 32'd0;
               A_SINT_CC_MAPR10NoCE1_ARA0_AD0 = 13'd0;
               end 
              if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==2'd2/*MS*/) && (xpc10nz==10'd540/*US*/) && !xpc10_stall)  begin 
               A_SINT_CC_MAPR10NoCE2_ARA0_WRD0 = 32'd0;
               A_SINT_CC_MAPR10NoCE2_ARA0_AD0 = 13'd0;
               end 
              if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==0/*MS*/) && (xpc10nz==10'd544/*US*/) && !xpc10_stall)  begin 
               A_SINT_CC_MAPR10NoCE0_ARA0_WRD0 = 32'd0;
               A_SINT_CC_MAPR10NoCE0_ARA0_AD0 = 13'd0;
               end 
              if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==1'd1/*MS*/) && (xpc10nz==10'd544/*US*/) && !xpc10_stall)  begin 
               A_SINT_CC_MAPR10NoCE1_ARA0_WRD0 = 32'd0;
               A_SINT_CC_MAPR10NoCE1_ARA0_AD0 = 13'd0;
               end 
              if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==0/*MS*/) && (xpc10nz==10'd547/*US*/) && !xpc10_stall)  begin 
               A_SINT_CC_MAPR10NoCE0_ARA0_WRD0 = 32'd0;
               A_SINT_CC_MAPR10NoCE0_ARA0_AD0 = 13'd0;
               end 
              
      case (xpc10nz) // synthesis full_case 
          10'd550/*US*/:  begin 
              if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==0/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE0_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE0_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==1'd1/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE1_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE1_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==2'd2/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE2_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE2_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==2'd3/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE3_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE3_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==0/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE0_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE0_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==1'd1/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE1_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE1_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==2'd2/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE2_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE2_ARA0_AD0 = 13'd0;
                       end 
                       end 
              
          10'd558/*US*/:  begin 
              if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [2'd3]==0/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE0_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE0_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [2'd3]==1'd1/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE1_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE1_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [2'd3]==2'd2/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE2_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE2_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [2'd3]==2'd3/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE3_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE3_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==0/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE0_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE0_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==1'd1/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE1_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE1_ARA0_AD0 = 13'd0;
                       end 
                       end 
              
          10'd565/*US*/:  begin 
              if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==0/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE0_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE0_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==1'd1/*MS*/) && !xpc10_stall
              )  begin 
                       A_SINT_CC_MAPR10NoCE1_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE1_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==2'd2/*MS*/) && !xpc10_stall
              )  begin 
                       A_SINT_CC_MAPR10NoCE2_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE2_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==2'd3/*MS*/) && !xpc10_stall
              )  begin 
                       A_SINT_CC_MAPR10NoCE3_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE3_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==0/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE0_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE0_ARA0_AD0 = 13'd0;
                       end 
                       end 
              endcase
      if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==0/*MS*/) && (xpc10nz==10'd571/*US*/) && !xpc10_stall)  begin 
               A_SINT_CC_MAPR10NoCE0_ARA0_WRD0 = 32'd0;
               A_SINT_CC_MAPR10NoCE0_ARA0_AD0 = 13'd0;
               end 
              
      case (xpc10nz) // synthesis full_case 
          10'd571/*US*/:  begin 
              if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==1'd1/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE1_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE1_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==2'd2/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE2_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE2_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==2'd3/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE3_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE3_ARA0_AD0 = 13'd0;
                       end 
                       end 
              
          10'd576/*US*/:  begin 
              if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [2'd3]==0/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE0_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE0_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [2'd3]==1'd1/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE1_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE1_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [2'd3]==2'd2/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE2_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE2_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [2'd3]==2'd3/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE3_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE3_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==0/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE0_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE0_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==1'd1/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE1_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE1_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==2'd2/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE2_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE2_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==2'd3/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE3_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE3_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]==0/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE0_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE0_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]==1'd1/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE1_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE1_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]==2'd2/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE2_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE2_ARA0_AD0 = 13'd0;
                       end 
                       end 
              
          10'd588/*US*/:  begin 
              if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==0/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE0_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE0_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==1'd1/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE1_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE1_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==2'd2/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE2_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE2_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==2'd3/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE3_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE3_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [2'd2]==0/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE0_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE0_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [2'd2]==1'd1/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE1_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE1_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [2'd2]==2'd2/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE2_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE2_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [2'd2]==2'd3/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE3_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE3_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]==0/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE0_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE0_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]==1'd1/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE1_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE1_ARA0_AD0 = 13'd0;
                       end 
                       end 
              
          10'd599/*US*/:  begin 
              if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==0/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE0_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE0_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==1'd1/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE1_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE1_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==2'd2/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE2_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE2_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && 
              (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==2'd3/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE3_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE3_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==0/*MS*/) && !xpc10_stall) 
               begin 
                       A_SINT_CC_MAPR10NoCE0_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE0_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==1'd1/*MS*/) && !xpc10_stall
              )  begin 
                       A_SINT_CC_MAPR10NoCE1_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE1_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==2'd2/*MS*/) && !xpc10_stall
              )  begin 
                       A_SINT_CC_MAPR10NoCE2_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE2_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==2'd3/*MS*/) && !xpc10_stall
              )  begin 
                       A_SINT_CC_MAPR10NoCE3_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE3_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]==0/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE0_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE0_ARA0_AD0 = 13'd0;
                       end 
                       end 
              
          10'd609/*US*/:  begin 
              if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==0/*MS*/) && !xpc10_stall
              )  begin 
                       A_SINT_CC_MAPR10NoCE0_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE0_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==1'd1/*MS*/) && 
              !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE1_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE1_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==2'd2/*MS*/) && 
              !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE2_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE2_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
              [2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==2'd3/*MS*/) && 
              !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE3_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE3_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==0/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE0_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE0_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==1'd1/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE1_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE1_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==2'd2/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE2_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE2_ARA0_AD0 = 13'd0;
                       end 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==2'd3/*MS*/) && !xpc10_stall)  begin 
                       A_SINT_CC_MAPR10NoCE3_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_MAPR10NoCE3_ARA0_AD0 = 13'd0;
                       end 
                       end 
              endcase
      if ((TTMT4Main_V_4>=15'h_5555) && !xpc10_stall)  begin if ((xpc10nz==8'd253/*US*/))  KppWaypoint0 = "Data Entered";
               end 
          if ((xpc10nz==7'd99/*US*/))  begin if ((TTMT4Main_V_10>=15'h_5555) && !xpc10_stall)  KppWaypoint0 = "Readback Done";
               end 
          if ((TTMT4Main_V_4>=15'h_5555) && !xpc10_stall)  begin if ((xpc10nz==7'd86/*US*/))  KppWaypoint0 = "Data Entered";
               end 
          if ((xpc10nz==7'd65/*US*/))  begin if ((TCCl0_12_V_0>=A_SINT_CC_SCALbx24_waycap) && !xpc10_stall)  KppWaypoint0 = "Cache Cleared"
              ;

               end 
          if (!xpc10_stall)  begin if ((xpc10nz==1'd1/*US*/))  KppWaypoint0 = "Start";
               end 
           end 
      

 always   @(posedge clk )  begin 
      //Start structure HPR cuckoo_hash_demo.exe
      if (reset)  begin 
               TCha6_10_V_0 <= 32'd0;
               A_SINT_CC_SCALbx24_next_victim <= 32'd0;
               fastspilldup26 <= 32'd0;
               TCin1_9_V_7 <= 32'd0;
               TCin1_9_V_6 <= 32'd0;
               A_SINT_CC_SCALbx24_stats_insert_evictions <= 32'd0;
               A_SINT_CC_SCALbx24_stats_insert_probes <= 32'd0;
               TCin1_9_V_5 <= 32'd0;
               TCin1_9_V_4 <= 32'd0;
               A_SINT_CC_SCALbx24_stats_inserts <= 32'd0;
               TCin1_9_V_3 <= 32'd0;
               A_SINT_CC_SCALbx24_next_free <= 32'd0;
               TCi1_SPILL_256 <= 32'd0;
               TTMT4Main_V_7 <= 32'd0;
               fastspilldup16 <= 32'd0;
               TCin1_9_V_1 <= 32'd0;
               TCin1_9_V_2 <= 32'd0;
               TTMT4Main_V_6 <= 64'd0;
               TCin1_9_V_0 <= 32'd0;
               fastspilldup12 <= 64'd0;
               TDGe1_4_V_0 <= 64'd0;
               TTMT4Main_V_5 <= 32'd0;
               TClo6_9_V_2 <= 32'd0;
               TCha3_10_V_0 <= 32'd0;
               A_SINT_CC_SCALbx24_stats_lookup_probes <= 32'd0;
               TClo6_9_V_0 <= 32'd0;
               done <= 1'd0;
               TTMT4Main_V_14 <= 32'd0;
               TCl6_SPILL_256 <= 32'd0;
               TClo6_9_V_1 <= 32'd0;
               TTMT4Main_V_13 <= 64'd0;
               A_SINT_CC_SCALbx24_stats_lookups <= 32'd0;
               TTMT4Main_V_12 <= 64'd0;
               fastspilldup30 <= 64'd0;
               TDGe6_4_V_0 <= 64'd0;
               TTMT4Main_V_11 <= 32'd0;
               TTMT4Main_V_10 <= 32'd0;
               TTMT4Main_V_8 <= 32'd0;
               TTMT4Main_V_9 <= 32'd0;
               TTMT4Main_V_3 <= 32'd0;
               TTMT4Main_V_4 <= 32'd0;
               TTMT4Main_V_2 <= 32'd0;
               A_SINT_CC_SCALbx28_seed <= 32'd0;
               A_64_US_CC_SCALbx28_dk <= 64'd0;
               TCCl0_12_V_0 <= 32'd0;
               TCCl0_12_V_1 <= 32'd0;
               A_SINT_CC_SCALbx24_waycap <= 32'd0;
               Z64USCCSCALbx26ARA0RRh10hold <= 64'd0;
               SINTCCMAPR12NoCE3ARB0RRh10hold <= 32'd0;
               SINTCCMAPR12NoCE2ARB0RRh10hold <= 32'd0;
               SINTCCMAPR12NoCE1ARB0RRh10hold <= 32'd0;
               SINTCCMAPR12NoCE0ARB0RRh10hold <= 32'd0;
               isMODULUS10RRh10primed <= 1'd0;
               isMODULUS10RRh10vld <= 1'd0;
               isMODULUS10RRh10hold <= 32'd0;
               SINTCCMAPR10NoCE3ARA0RRh10hold <= 32'd0;
               SINTCCMAPR10NoCE2ARA0RRh10hold <= 32'd0;
               SINTCCMAPR10NoCE1ARA0RRh10hold <= 32'd0;
               SINTCCMAPR10NoCE0ARA0RRh10hold <= 32'd0;
               SINTCCMAPR10NoCE0ARA0RRh10shot0 <= 1'd0;
               SINTCCMAPR10NoCE1ARA0RRh10shot0 <= 1'd0;
               SINTCCMAPR10NoCE2ARA0RRh10shot0 <= 1'd0;
               SINTCCMAPR10NoCE3ARA0RRh10shot0 <= 1'd0;
               SINTCCMAPR12NoCE0ARB0RRh10shot0 <= 1'd0;
               SINTCCMAPR12NoCE1ARB0RRh10shot0 <= 1'd0;
               SINTCCMAPR12NoCE2ARB0RRh10shot0 <= 1'd0;
               SINTCCMAPR12NoCE3ARB0RRh10shot0 <= 1'd0;
               Z64USCCSCALbx26ARA0RRh10shot0 <= 1'd0;
               xpc10_trk64 <= 1'd0;
               xpc10_trk63 <= 1'd0;
               xpc10_trk62 <= 1'd0;
               xpc10_trk61 <= 1'd0;
               xpc10_trk60 <= 1'd0;
               xpc10_trk59 <= 1'd0;
               xpc10_trk58 <= 1'd0;
               xpc10_trk57 <= 1'd0;
               xpc10_trk56 <= 1'd0;
               xpc10_trk55 <= 1'd0;
               xpc10_trk54 <= 1'd0;
               xpc10_trk53 <= 1'd0;
               xpc10_trk52 <= 1'd0;
               xpc10_trk51 <= 1'd0;
               xpc10_trk50 <= 1'd0;
               xpc10_trk49 <= 1'd0;
               xpc10_trk48 <= 1'd0;
               xpc10_trk47 <= 1'd0;
               xpc10_trk46 <= 1'd0;
               xpc10_trk45 <= 1'd0;
               xpc10_trk44 <= 1'd0;
               xpc10_trk43 <= 1'd0;
               xpc10_trk42 <= 1'd0;
               xpc10_trk41 <= 1'd0;
               xpc10_trk40 <= 1'd0;
               xpc10_trk39 <= 1'd0;
               xpc10_trk38 <= 1'd0;
               xpc10_trk37 <= 1'd0;
               xpc10_trk36 <= 1'd0;
               xpc10_trk35 <= 1'd0;
               xpc10_trk34 <= 1'd0;
               xpc10_trk33 <= 1'd0;
               xpc10_trk32 <= 1'd0;
               xpc10_trk31 <= 1'd0;
               xpc10_trk30 <= 1'd0;
               xpc10_trk29 <= 1'd0;
               xpc10_trk28 <= 1'd0;
               xpc10_trk27 <= 1'd0;
               xpc10_trk26 <= 1'd0;
               xpc10_trk25 <= 1'd0;
               xpc10_trk24 <= 1'd0;
               xpc10_trk23 <= 1'd0;
               xpc10_trk22 <= 1'd0;
               xpc10_trk21 <= 1'd0;
               xpc10_trk20 <= 1'd0;
               xpc10_trk19 <= 1'd0;
               xpc10_trk18 <= 1'd0;
               xpc10_trk17 <= 1'd0;
               xpc10_trk16 <= 1'd0;
               xpc10_trk15 <= 1'd0;
               xpc10_trk14 <= 1'd0;
               xpc10_trk13 <= 1'd0;
               xpc10_trk12 <= 1'd0;
               xpc10_trk11 <= 1'd0;
               xpc10_trk10 <= 1'd0;
               xpc10_trk9 <= 1'd0;
               xpc10_trk8 <= 1'd0;
               xpc10_trk7 <= 1'd0;
               xpc10_trk6 <= 1'd0;
               xpc10_trk5 <= 1'd0;
               xpc10_trk4 <= 1'd0;
               xpc10_trk3 <= 1'd0;
               xpc10_trk2 <= 1'd0;
               xpc10_trk1 <= 1'd0;
               xpc10_trk0 <= 1'd0;
               xpc10nz <= 10'd0;
               end 
               else  begin 
              if ((!xpc10_stall || (TCin1_9_V_4<3'd4)) && (xpc10nz==9'd503/*US*/) && (TCin1_9_V_4==3'd4/*US*/)) $display("Eviction %1d needed"
                  , TCin1_9_V_1);
                  if ((xpc10nz==9'd473/*US*/))  begin 
                      if (((xpc10nz==9'd473/*US*/)? !A_SINT_CC_MAPR10NoCE3_ARA0_RDD0 && !xpc10_stall: !SINTCCMAPR10NoCE3ARA0RRh10hold
                       && !xpc10_stall) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd3/*MS*/) && (TCin1_9_V_4==3'd4/*US*/)) $display("Eviction %1d needed"
                          , TCin1_9_V_1);
                          if (((xpc10nz==9'd473/*US*/)? !A_SINT_CC_MAPR10NoCE2_ARA0_RDD0 && !xpc10_stall: !SINTCCMAPR10NoCE2ARA0RRh10hold
                       && !xpc10_stall) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd2/*MS*/) && (TCin1_9_V_4==3'd4/*US*/)) $display("Eviction %1d needed"
                          , TCin1_9_V_1);
                          if (((xpc10nz==9'd473/*US*/)? !A_SINT_CC_MAPR10NoCE1_ARA0_RDD0 && !xpc10_stall: !SINTCCMAPR10NoCE1ARA0RRh10hold
                       && !xpc10_stall) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==1'd1/*MS*/) && (TCin1_9_V_4==3'd4/*US*/)) $display("Eviction %1d needed"
                          , TCin1_9_V_1);
                          if (((xpc10nz==9'd473/*US*/)? !A_SINT_CC_MAPR10NoCE0_ARA0_RDD0 && !xpc10_stall: !SINTCCMAPR10NoCE0ARA0RRh10hold
                       && !xpc10_stall) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==0/*MS*/) && (TCin1_9_V_4==3'd4/*US*/)) $display("Eviction %1d needed"
                          , TCin1_9_V_1);
                          if ((TCin1_9_V_4==3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [TCin1_9_V_4]!=0/*MS*/) && !xpc10_stall) $display("Eviction %1d needed", TCin1_9_V_1);
                           end 
                      if ((!xpc10_stall || (TCin1_9_V_4<3'd4)) && (xpc10nz==9'd259/*US*/) && (TCin1_9_V_4==3'd4/*US*/)) $display("Eviction %1d needed"
                  , TCin1_9_V_1);
                  if ((TTMT4Main_V_4>=15'h_5555) && (xpc10nz==8'd253/*US*/) && !xpc10_stall) $display("Cuckoo cache inserted items %1d/%1d"
                  , TTMT4Main_V_3, TTMT4Main_V_2);
                  if (!xpc10_stall) 
                  case (xpc10nz) // synthesis full_case 
                      7'd100/*US*/:  begin 
                          $display("cuckoo cache: this=%1d, inserts=%1d, lookups=%1d", 0, A_SINT_CC_SCALbx24_stats_inserts, A_SINT_CC_SCALbx24_stats_lookups
                          );
                          $display("cuckoo cache: insert_probes=%1d, insert_evictions=%1d", A_SINT_CC_SCALbx24_stats_insert_probes, A_SINT_CC_SCALbx24_stats_insert_evictions
                          );
                           end 
                          
                      7'd101/*US*/:  begin 
                          $display("cuckoo cache: lookup_probes=%1d", A_SINT_CC_SCALbx24_stats_lookup_probes);
                          $display("Cuckoo cache demo finished.");
                           end 
                          
                      7'd102/*US*/: $finish(0);
                  endcase
                  if ((xpc10nz==7'd99/*US*/))  begin if ((TTMT4Main_V_10>=15'h_5555) && !xpc10_stall) $display("Cuckoo cache inserted items %1d/%1d"
                      , TTMT4Main_V_9, TTMT4Main_V_8);
                       end 
                  if ((TTMT4Main_V_4>=15'h_5555) && (xpc10nz==7'd86/*US*/) && !xpc10_stall) $display("Cuckoo cache inserted items %1d/%1d"
                  , TTMT4Main_V_3, TTMT4Main_V_2);
                  if ((xpc10nz==7'd65/*US*/))  begin if ((TCCl0_12_V_0>=A_SINT_CC_SCALbx24_waycap) && !xpc10_stall) $display("Cuckoo cache cleared"
                      );
                       end 
                  if (!xpc10_stall) 
                  case (xpc10nz) // synthesis full_case 
                      1'd1/*US*/: $display("Cuckoo cache testbench start. Capacity=%1d", 16'h_8000);

                      3'd4/*US*/:  A_SINT_CC_SCALbx24_waycap <= 32'h_2000;

                      3'd5/*US*/:  A_sA_SINT_CC_SCALbx20_ARA0[0] <= 32'd0;

                      3'd7/*US*/:  A_sA_SINT_CC_SCALbx20_ARA0[1'd1] <= 32'd1;

                      4'd8/*US*/:  A_sA_SINT_CC_SCALbx20_ARA0[2'd2] <= 32'd2;

                      4'd10/*US*/:  A_sA_SINT_CC_SCALbx20_ARA0[2'd3] <= 32'd3;

                      4'd12/*US*/:  A_sA_SINT_CC_SCALbx22_ARB0[0] <= 32'd0;

                      4'd13/*US*/:  A_sA_SINT_CC_SCALbx22_ARB0[1'd1] <= 32'd1;

                      4'd15/*US*/:  A_sA_SINT_CC_SCALbx22_ARB0[2'd2] <= 32'd2;

                      5'd16/*US*/:  A_sA_SINT_CC_SCALbx22_ARB0[2'd3] <= 32'd3;

                      5'd19/*US*/:  begin 
                           TCCl0_12_V_0 <= 32'd0;
                           TCCl0_12_V_1 <= 32'd0;
                           end 
                          
                      7'd64/*US*/:  TCCl0_12_V_0 <= 32'd1+TCCl0_12_V_0;

                      7'd82/*US*/:  begin 
                           A_SINT_CC_SCALbx28_seed <= 32'h1_e240;
                           A_64_US_CC_SCALbx28_dk <= 64'h23_86f2_69cb_1f00;
                           end 
                          
                      7'd83/*US*/:  A_SINT_CC_SCALbx28_seed <= 32'h1_e240;

                      7'd84/*US*/:  begin 
                           TTMT4Main_V_2 <= 32'd0;
                           A_64_US_CC_SCALbx28_dk <= 64'h23_86f2_69cb_1f00;
                           end 
                          
                      7'd85/*US*/:  begin 
                           TTMT4Main_V_3 <= 32'd0;
                           TTMT4Main_V_4 <= 32'd0;
                           end 
                          
                      7'd87/*US*/:  begin 
                           A_SINT_CC_SCALbx28_seed <= 32'h1_e240;
                           A_64_US_CC_SCALbx28_dk <= 64'h23_86f2_69cb_1f00;
                           end 
                          
                      7'd88/*US*/:  begin 
                           TTMT4Main_V_8 <= 32'd0;
                           TTMT4Main_V_9 <= 32'd0;
                           end 
                          
                      7'd89/*US*/:  begin 
                           TTMT4Main_V_10 <= 32'd0;
                           A_SINT_CC_SCALbx28_seed <= 32'h_2aa0_1d31+32'h_7ff8_a3ed*A_SINT_CC_SCALbx28_seed;
                           end 
                          
                      7'd90/*US*/:  TTMT4Main_V_11 <= A_SINT_CC_SCALbx28_seed;

                      7'd91/*US*/:  begin 
                           fastspilldup30 <= A_64_US_CC_SCALbx28_dk;
                           TDGe6_4_V_0 <= A_64_US_CC_SCALbx28_dk;
                           end 
                          
                      7'd92/*US*/:  A_64_US_CC_SCALbx28_dk <= 64'h1+fastspilldup30;

                      7'd93/*US*/:  TTMT4Main_V_12 <= TDGe6_4_V_0;

                      7'd94/*US*/:  A_SINT_CC_SCALbx24_stats_lookups <= 32'd1+A_SINT_CC_SCALbx24_stats_lookups;

                      7'd97/*US*/:  TTMT4Main_V_8 <= 32'd1+TTMT4Main_V_8;

                      7'd98/*US*/:  TTMT4Main_V_10 <= 32'd1+TTMT4Main_V_10;

                      7'd102/*US*/:  done <= 1'h1;

                      7'd103/*US*/:  TClo6_9_V_0 <= 32'd0;

                      7'd104/*US*/:  A_SINT_CC_SCALbx24_stats_lookup_probes <= 32'd1+A_SINT_CC_SCALbx24_stats_lookup_probes;

                      7'd105/*US*/:  TCha3_10_V_0 <= TTMT4Main_V_11+32'd51*TClo6_9_V_0;

                      8'd235/*US*/:  TClo6_9_V_1 <= (isMODULUS10RRh10vld? isMODULUS10RRh10hold: isMODULUS10_RR);

                      8'd240/*US*/:  TTMT4Main_V_13 <= ((xpc10nz==8'd240/*US*/)? A_64_US_CC_SCALbx26_ARA0_RDD0: Z64USCCSCALbx26ARA0RRh10hold
                      );


                      8'd241/*US*/:  begin 
                           TTMT4Main_V_14 <= 32'h0;
                           TCl6_SPILL_256 <= 32'd0;
                           end 
                          
                      8'd244/*US*/:  TTMT4Main_V_5 <= A_SINT_CC_SCALbx28_seed;

                      8'd245/*US*/:  begin 
                           fastspilldup12 <= A_64_US_CC_SCALbx28_dk;
                           TDGe1_4_V_0 <= A_64_US_CC_SCALbx28_dk;
                           end 
                          
                      8'd246/*US*/:  A_64_US_CC_SCALbx28_dk <= 64'h1+fastspilldup12;

                      8'd247/*US*/:  begin 
                           TTMT4Main_V_6 <= TDGe1_4_V_0;
                           TCin1_9_V_0 <= TTMT4Main_V_5;
                           end 
                          
                      8'd248/*US*/:  begin 
                           TCin1_9_V_1 <= 32'd0;
                           TCin1_9_V_2 <= 32'd0;
                           end 
                          
                      8'd251/*US*/:  TTMT4Main_V_2 <= 32'd1+TTMT4Main_V_2;

                      8'd252/*US*/:  TTMT4Main_V_4 <= 32'd1+TTMT4Main_V_4;

                      8'd254/*US*/:  begin 
                           TCin1_9_V_3 <= fastspilldup16;
                           A_SINT_CC_SCALbx24_next_free <= 32'd1+fastspilldup16;
                           end 
                          
                      8'd255/*US*/:  TCin1_9_V_2 <= TCin1_9_V_3;

                      9'd257/*US*/:  A_SINT_CC_SCALbx24_stats_inserts <= 32'd1+A_SINT_CC_SCALbx24_stats_inserts;

                      9'd258/*US*/:  begin 
                           TCin1_9_V_5 <= 32'd0;
                           TCin1_9_V_4 <= 32'd0;
                           end 
                          
                      9'd284/*US*/:  A_SINT_CC_SCALbx24_stats_insert_evictions <= 32'd1+A_SINT_CC_SCALbx24_stats_insert_evictions;

                      9'd286/*US*/:  TCin1_9_V_6 <= ((A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]==2'd3/*MS*/)? ((xpc10nz
                      ==9'd286/*US*/)? A_SINT_CC_MAPR10NoCE3_ARA0_RDD0: SINTCCMAPR10NoCE3ARA0RRh10hold): ((A_sA_SINT_CC_SCALbx20_ARA0
                      [A_SINT_CC_SCALbx24_next_victim]==2'd2/*MS*/)? ((xpc10nz==9'd286/*US*/)? A_SINT_CC_MAPR10NoCE2_ARA0_RDD0: SINTCCMAPR10NoCE2ARA0RRh10hold
                      ): ((A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]==1'd1/*MS*/)? ((xpc10nz==9'd286/*US*/)? A_SINT_CC_MAPR10NoCE1_ARA0_RDD0
                      : SINTCCMAPR10NoCE1ARA0RRh10hold): ((A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]==0/*MS*/)? ((xpc10nz
                      ==9'd286/*US*/)? A_SINT_CC_MAPR10NoCE0_ARA0_RDD0: SINTCCMAPR10NoCE0ARA0RRh10hold): 32'bx))));


                      9'd288/*US*/:  TCin1_9_V_7 <= ((A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]==2'd3/*MS*/)? ((xpc10nz
                      ==9'd288/*US*/)? A_SINT_CC_MAPR12NoCE3_ARB0_RDD0: SINTCCMAPR12NoCE3ARB0RRh10hold): ((A_sA_SINT_CC_SCALbx22_ARB0
                      [A_SINT_CC_SCALbx24_next_victim]==2'd2/*MS*/)? ((xpc10nz==9'd288/*US*/)? A_SINT_CC_MAPR12NoCE2_ARB0_RDD0: SINTCCMAPR12NoCE2ARB0RRh10hold
                      ): ((A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]==1'd1/*MS*/)? ((xpc10nz==9'd288/*US*/)? A_SINT_CC_MAPR12NoCE1_ARB0_RDD0
                      : SINTCCMAPR12NoCE1ARB0RRh10hold): ((A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]==0/*MS*/)? ((xpc10nz
                      ==9'd288/*US*/)? A_SINT_CC_MAPR12NoCE0_ARB0_RDD0: SINTCCMAPR12NoCE0ARB0RRh10hold): 32'bx))));


                      9'd318/*US*/:  TCin1_9_V_2 <= TCin1_9_V_7;

                      9'd319/*US*/:  fastspilldup26 <= 32'd1+A_SINT_CC_SCALbx24_next_victim;

                      9'd320/*US*/:  begin 
                           A_SINT_CC_SCALbx24_next_victim <= fastspilldup26;
                           TCin1_9_V_3 <= fastspilldup26;
                           end 
                          
                      9'd321/*US*/:  A_SINT_CC_SCALbx24_next_victim <= (TCin1_9_V_3%3'd4);

                      9'd322/*US*/:  begin 
                           TCin1_9_V_5 <= 32'd0;
                           TCin1_9_V_4 <= 32'd0;
                           end 
                          
                      9'd323/*US*/:  fastspilldup26 <= 32'd1+A_SINT_CC_SCALbx24_next_victim;

                      9'd329/*US*/:  begin 
                           TCin1_9_V_2 <= TCin1_9_V_7;
                           TCin1_9_V_0 <= TCin1_9_V_6;
                           end 
                          
                      9'd340/*US*/:  begin 
                           TCi1_SPILL_256 <= 32'd0;
                           TTMT4Main_V_7 <= 32'h0;
                           end 
                          
                      9'd341/*US*/:  TCha6_10_V_0 <= TCin1_9_V_0+32'd51*TCin1_9_V_4;

                      9'd471/*US*/:  TCin1_9_V_5 <= (isMODULUS10RRh10vld? isMODULUS10RRh10hold: isMODULUS10_RR);

                      9'd502/*US*/:  TCin1_9_V_1 <= 32'd1+TCin1_9_V_1;

                      10'd537/*US*/:  TCCl0_12_V_1 <= 32'd1+TCCl0_12_V_1;

                      10'd539/*US*/:  TCCl0_12_V_1 <= 32'd1+TCCl0_12_V_1;

                      10'd549/*US*/:  begin 
                           TCCl0_12_V_0 <= 32'd1+TCCl0_12_V_0;
                           TCCl0_12_V_1 <= 32'd4;
                           end 
                          endcase
                  
              case (xpc10nz) // synthesis full_case 
                  5'd20/*US*/:  begin 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd3]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=1'd1
                      /*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=0/*MS*/) && !xpc10_stall)  begin 
                               TCCl0_12_V_0 <= 32'd1+TCCl0_12_V_0;
                               TCCl0_12_V_1 <= 32'd4;
                               end 
                              if ((A_sA_SINT_CC_SCALbx20_ARA0[0]==2'd3/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd1;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[0]==2'd2/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd1;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[0]==1'd1/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd1;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[0]==0/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd1;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]==2'd3/*MS*/) && 
                      !xpc10_stall)  TCCl0_12_V_1 <= 32'd1;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]==2'd2/*MS*/) && 
                      !xpc10_stall)  TCCl0_12_V_1 <= 32'd1;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]==1'd1/*MS*/) && 
                      !xpc10_stall)  TCCl0_12_V_1 <= 32'd1;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]==0/*MS*/) && 
                      !xpc10_stall)  TCCl0_12_V_1 <= 32'd1;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==2'd3/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd2;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==2'd2/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd2;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==1'd1/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd2;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==0/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd2;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd3]==2'd3/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd3;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd3]==2'd2/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd3;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd3]==1'd1/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd3;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd3]==0/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd3;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[0]==2'd3/*MS*/))  xpc10nz <= 5'd21/*US*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[0]==2'd2/*MS*/))  xpc10nz <= 5'd22/*US*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[0]==1'd1/*MS*/))  xpc10nz <= 5'd23/*US*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[0]==0/*MS*/))  xpc10nz <= 5'd24/*US*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]==2'd3/*MS*/)) 
                       xpc10nz <= 5'd25/*US*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]==2'd2/*MS*/)) 
                       xpc10nz <= 5'd26/*US*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]==1'd1/*MS*/)) 
                       xpc10nz <= 5'd27/*US*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]==0/*MS*/))  xpc10nz
                           <= 5'd28/*US*/;

                          if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==2'd3/*MS*/))  xpc10nz <= 5'd29/*US*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==2'd2/*MS*/))  xpc10nz <= 5'd30/*US*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==1'd1/*MS*/))  xpc10nz <= 5'd31/*US*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==0/*MS*/))  xpc10nz <= 6'd32/*US*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd3]==2'd3/*MS*/))  xpc10nz <= 6'd33/*US*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd3]==2'd2/*MS*/))  xpc10nz <= 6'd34/*US*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd3]==1'd1/*MS*/))  xpc10nz <= 6'd35/*US*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd3]==0/*MS*/))  xpc10nz <= 6'd36/*US*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd3]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=1'd1
                      /*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=0/*MS*/))  xpc10nz <= 7'd65/*xpc10nz*/;
                           end 
                      
                  6'd37/*US*/:  begin 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]==0/*MS*/))  xpc10nz <= 6'd41/*US*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]==0/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd2;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]==1'd1/*MS*/))  xpc10nz <= 6'd40/*US*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]==1'd1/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd2;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]==2'd2/*MS*/))  xpc10nz <= 6'd39/*US*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=2'd2/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=0/*MS*/) && !xpc10_stall) 
                       begin 
                               TCCl0_12_V_0 <= 32'd1+TCCl0_12_V_0;
                               TCCl0_12_V_1 <= 32'd4;
                               end 
                              if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]==2'd2/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd2;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]==2'd3/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd2;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==2'd3/*MS*/) && 
                      !xpc10_stall)  TCCl0_12_V_1 <= 32'd2;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==2'd2/*MS*/) && 
                      !xpc10_stall)  TCCl0_12_V_1 <= 32'd2;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==1'd1/*MS*/) && 
                      !xpc10_stall)  TCCl0_12_V_1 <= 32'd2;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==0/*MS*/) && 
                      !xpc10_stall)  TCCl0_12_V_1 <= 32'd2;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==2'd3/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd3;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==2'd2/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd3;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==1'd1/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd3;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==0/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd3;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]==2'd3/*MS*/))  xpc10nz <= 6'd38/*US*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==2'd3/*MS*/)) 
                       xpc10nz <= 6'd42/*US*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==2'd2/*MS*/)) 
                       xpc10nz <= 6'd43/*US*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==1'd1/*MS*/)) 
                       xpc10nz <= 6'd44/*US*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==0/*MS*/)) 
                       xpc10nz <= 6'd45/*US*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==2'd3/*MS*/))  xpc10nz <= 6'd46/*US*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==2'd2/*MS*/))  xpc10nz <= 6'd47/*US*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==1'd1/*MS*/))  xpc10nz <= 6'd48/*US*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==0/*MS*/))  xpc10nz <= 6'd49/*US*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=2'd2/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=0/*MS*/))  xpc10nz <= 7'd65
                          /*xpc10nz*/;

                           end 
                      
                  6'd50/*US*/:  begin 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==0/*MS*/))  xpc10nz <= 6'd54/*US*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==0/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd3;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==1'd1/*MS*/))  xpc10nz <= 6'd53/*US*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd3]!=0/*MS*/) && !xpc10_stall)  begin 
                               TCCl0_12_V_0 <= 32'd1+TCCl0_12_V_0;
                               TCCl0_12_V_1 <= 32'd4;
                               end 
                              if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==1'd1/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd3;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==2'd2/*MS*/))  xpc10nz <= 6'd52/*US*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==2'd2/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd3;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd3]!=0/*MS*/))  xpc10nz <= 7'd65/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==0/*MS*/)) 
                       xpc10nz <= 6'd58/*US*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==1'd1/*MS*/)) 
                       xpc10nz <= 6'd57/*US*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==2'd2/*MS*/)) 
                       xpc10nz <= 6'd56/*US*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==2'd3/*MS*/)) 
                       xpc10nz <= 6'd55/*US*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==2'd3/*MS*/))  xpc10nz <= 6'd51/*US*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==0/*MS*/) && 
                      !xpc10_stall)  TCCl0_12_V_1 <= 32'd3;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==1'd1/*MS*/) && 
                      !xpc10_stall)  TCCl0_12_V_1 <= 32'd3;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==2'd2/*MS*/) && 
                      !xpc10_stall)  TCCl0_12_V_1 <= 32'd3;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==2'd3/*MS*/) && 
                      !xpc10_stall)  TCCl0_12_V_1 <= 32'd3;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==2'd3/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd3;
                           end 
                      
                  6'd59/*US*/:  begin 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==0/*MS*/))  xpc10nz <= 6'd63/*US*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==0/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd4;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==1'd1/*MS*/))  xpc10nz <= 6'd62/*US*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd3]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=0/*MS*/) && !xpc10_stall)  begin 
                               TCCl0_12_V_0 <= 32'd1+TCCl0_12_V_0;
                               TCCl0_12_V_1 <= 32'd4;
                               end 
                              if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==1'd1/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd4;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==2'd2/*MS*/))  xpc10nz <= 6'd61/*US*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==2'd2/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd4;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd3]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=0/*MS*/))  xpc10nz <= 7'd65/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==2'd3/*MS*/))  xpc10nz <= 6'd60/*US*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==2'd3/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd4;
                           end 
                      
                  7'd65/*US*/:  begin 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd3]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=1'd1
                      /*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=0/*MS*/) && (TCCl0_12_V_0<A_SINT_CC_SCALbx24_waycap) && !xpc10_stall
                      )  begin 
                               TCCl0_12_V_0 <= 32'd1+TCCl0_12_V_0;
                               TCCl0_12_V_1 <= 32'd4;
                               end 
                              if ((A_sA_SINT_CC_SCALbx20_ARA0[0]==2'd3/*MS*/) && (TCCl0_12_V_0<A_SINT_CC_SCALbx24_waycap) && !xpc10_stall
                      )  TCCl0_12_V_1 <= 32'd0;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[0]==2'd2/*MS*/) && (TCCl0_12_V_0<A_SINT_CC_SCALbx24_waycap) && !xpc10_stall
                      )  TCCl0_12_V_1 <= 32'd0;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[0]==1'd1/*MS*/) && (TCCl0_12_V_0<A_SINT_CC_SCALbx24_waycap) && !xpc10_stall
                      )  TCCl0_12_V_1 <= 32'd0;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[0]==0/*MS*/) && (TCCl0_12_V_0<A_SINT_CC_SCALbx24_waycap) && !xpc10_stall)  TCCl0_12_V_1
                           <= 32'd0;

                          if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]==2'd3/*MS*/) && 
                      (TCCl0_12_V_0<A_SINT_CC_SCALbx24_waycap) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd1;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]==2'd2/*MS*/) && 
                      (TCCl0_12_V_0<A_SINT_CC_SCALbx24_waycap) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd1;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]==1'd1/*MS*/) && 
                      (TCCl0_12_V_0<A_SINT_CC_SCALbx24_waycap) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd1;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]==0/*MS*/) && 
                      (TCCl0_12_V_0<A_SINT_CC_SCALbx24_waycap) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd1;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==2'd3/*MS*/) && (TCCl0_12_V_0<A_SINT_CC_SCALbx24_waycap) && 
                      !xpc10_stall)  TCCl0_12_V_1 <= 32'd2;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==2'd2/*MS*/) && (TCCl0_12_V_0<A_SINT_CC_SCALbx24_waycap) && 
                      !xpc10_stall)  TCCl0_12_V_1 <= 32'd2;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==1'd1/*MS*/) && (TCCl0_12_V_0<A_SINT_CC_SCALbx24_waycap) && 
                      !xpc10_stall)  TCCl0_12_V_1 <= 32'd2;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==0/*MS*/) && (TCCl0_12_V_0<A_SINT_CC_SCALbx24_waycap) && 
                      !xpc10_stall)  TCCl0_12_V_1 <= 32'd2;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd3]==2'd3/*MS*/) && (TCCl0_12_V_0<A_SINT_CC_SCALbx24_waycap) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd3;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd3]==2'd2/*MS*/) && (TCCl0_12_V_0<A_SINT_CC_SCALbx24_waycap) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd3;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd3]==1'd1/*MS*/) && (TCCl0_12_V_0<A_SINT_CC_SCALbx24_waycap) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd3;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd3]==0/*MS*/) && (TCCl0_12_V_0<A_SINT_CC_SCALbx24_waycap) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd3;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd3]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=1'd1
                      /*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=0/*MS*/) && (TCCl0_12_V_0<A_SINT_CC_SCALbx24_waycap))  xpc10nz <= 7'd65
                          /*xpc10nz*/;

                          if ((TCCl0_12_V_0>=A_SINT_CC_SCALbx24_waycap))  xpc10nz <= 7'd82/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[0]==2'd3/*MS*/) && (TCCl0_12_V_0<A_SINT_CC_SCALbx24_waycap))  xpc10nz <= 7'd66
                          /*xpc10nz*/;

                          if ((A_sA_SINT_CC_SCALbx20_ARA0[0]==2'd2/*MS*/) && (TCCl0_12_V_0<A_SINT_CC_SCALbx24_waycap))  xpc10nz <= 7'd67
                          /*xpc10nz*/;

                          if ((A_sA_SINT_CC_SCALbx20_ARA0[0]==1'd1/*MS*/) && (TCCl0_12_V_0<A_SINT_CC_SCALbx24_waycap))  xpc10nz <= 7'd68
                          /*xpc10nz*/;

                          if ((A_sA_SINT_CC_SCALbx20_ARA0[0]==0/*MS*/) && (TCCl0_12_V_0<A_SINT_CC_SCALbx24_waycap))  xpc10nz <= 7'd69
                          /*xpc10nz*/;

                          if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]==2'd3/*MS*/) && 
                      (TCCl0_12_V_0<A_SINT_CC_SCALbx24_waycap))  xpc10nz <= 7'd70/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]==2'd2/*MS*/) && 
                      (TCCl0_12_V_0<A_SINT_CC_SCALbx24_waycap))  xpc10nz <= 7'd71/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]==1'd1/*MS*/) && 
                      (TCCl0_12_V_0<A_SINT_CC_SCALbx24_waycap))  xpc10nz <= 7'd72/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]==0/*MS*/) && 
                      (TCCl0_12_V_0<A_SINT_CC_SCALbx24_waycap))  xpc10nz <= 7'd73/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==2'd3/*MS*/) && (TCCl0_12_V_0<A_SINT_CC_SCALbx24_waycap)) 
                       xpc10nz <= 7'd74/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==2'd2/*MS*/) && (TCCl0_12_V_0<A_SINT_CC_SCALbx24_waycap)) 
                       xpc10nz <= 7'd75/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==1'd1/*MS*/) && (TCCl0_12_V_0<A_SINT_CC_SCALbx24_waycap)) 
                       xpc10nz <= 7'd76/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==0/*MS*/) && (TCCl0_12_V_0<A_SINT_CC_SCALbx24_waycap))  xpc10nz
                           <= 7'd77/*xpc10nz*/;

                          if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd3]==2'd3/*MS*/) && (TCCl0_12_V_0<A_SINT_CC_SCALbx24_waycap))  xpc10nz <= 7'd78/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd3]==2'd2/*MS*/) && (TCCl0_12_V_0<A_SINT_CC_SCALbx24_waycap))  xpc10nz <= 7'd79/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd3]==1'd1/*MS*/) && (TCCl0_12_V_0<A_SINT_CC_SCALbx24_waycap))  xpc10nz <= 7'd80/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [0]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[0]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd3]==0/*MS*/) && (TCCl0_12_V_0<A_SINT_CC_SCALbx24_waycap))  xpc10nz <= 7'd81/*xpc10nz*/;
                           end 
                      
                  7'd96/*US*/:  begin 
                      if (!(!(32'hffffffff&TCl6_SPILL_256)) && !xpc10_stall)  begin 
                               TTMT4Main_V_14 <= TCl6_SPILL_256;
                               TTMT4Main_V_8 <= 32'd1+TTMT4Main_V_8;
                               end 
                              if ((TTMT4Main_V_12!=TTMT4Main_V_13) && !(32'hffffffff&TCl6_SPILL_256) && !xpc10_stall)  begin 
                               TTMT4Main_V_14 <= TCl6_SPILL_256;
                               TTMT4Main_V_8 <= 32'd1+TTMT4Main_V_8;
                               end 
                              if ((TTMT4Main_V_12==TTMT4Main_V_13) && !(32'hffffffff&TCl6_SPILL_256) && !xpc10_stall)  begin 
                               TTMT4Main_V_14 <= TCl6_SPILL_256;
                               TTMT4Main_V_9 <= 32'd1+TTMT4Main_V_9;
                               end 
                              if ((TTMT4Main_V_12==TTMT4Main_V_13) && !(32'hffffffff&TCl6_SPILL_256))  xpc10nz <= 7'd97/*xpc10nz*/;
                          if ((!(!(32'hffffffff&TCl6_SPILL_256))? 1'd1: (TTMT4Main_V_12!=TTMT4Main_V_13)))  xpc10nz <= 7'd98/*xpc10nz*/;
                           end 
                      
                  8'd237/*US*/:  begin 
                      if ((TClo6_9_V_0==3'd4/*US*/) && (TTMT4Main_V_11==((A_sA_SINT_CC_SCALbx20_ARA0[TClo6_9_V_0]==2'd3/*MS*/)? ((xpc10nz
                      ==8'd237/*US*/)? A_SINT_CC_MAPR10NoCE3_ARA0_RDD0: SINTCCMAPR10NoCE3ARA0RRh10hold): ((A_sA_SINT_CC_SCALbx20_ARA0
                      [TClo6_9_V_0]==2'd2/*MS*/)? ((xpc10nz==8'd237/*US*/)? A_SINT_CC_MAPR10NoCE2_ARA0_RDD0: SINTCCMAPR10NoCE2ARA0RRh10hold
                      ): ((A_sA_SINT_CC_SCALbx20_ARA0[TClo6_9_V_0]==1'd1/*MS*/)? ((xpc10nz==8'd237/*US*/)? A_SINT_CC_MAPR10NoCE1_ARA0_RDD0
                      : SINTCCMAPR10NoCE1ARA0RRh10hold): ((A_sA_SINT_CC_SCALbx20_ARA0[TClo6_9_V_0]==0/*MS*/)? ((xpc10nz==8'd237/*US*/)? A_SINT_CC_MAPR10NoCE0_ARA0_RDD0
                      : SINTCCMAPR10NoCE0ARA0RRh10hold): 1'bx))))) && !xpc10_stall)  begin 
                               TTMT4Main_V_14 <= -32'h5;
                               TCl6_SPILL_256 <= -32'd5;
                               end 
                              if ((TClo6_9_V_0!=3'd4/*US*/) && (TTMT4Main_V_11==((A_sA_SINT_CC_SCALbx20_ARA0[TClo6_9_V_0]==2'd3/*MS*/)? ((xpc10nz
                      ==8'd237/*US*/)? A_SINT_CC_MAPR10NoCE3_ARA0_RDD0: SINTCCMAPR10NoCE3ARA0RRh10hold): ((A_sA_SINT_CC_SCALbx20_ARA0
                      [TClo6_9_V_0]==2'd2/*MS*/)? ((xpc10nz==8'd237/*US*/)? A_SINT_CC_MAPR10NoCE2_ARA0_RDD0: SINTCCMAPR10NoCE2ARA0RRh10hold
                      ): ((A_sA_SINT_CC_SCALbx20_ARA0[TClo6_9_V_0]==1'd1/*MS*/)? ((xpc10nz==8'd237/*US*/)? A_SINT_CC_MAPR10NoCE1_ARA0_RDD0
                      : SINTCCMAPR10NoCE1ARA0RRh10hold): ((A_sA_SINT_CC_SCALbx20_ARA0[TClo6_9_V_0]==0/*MS*/)? ((xpc10nz==8'd237/*US*/)? A_SINT_CC_MAPR10NoCE0_ARA0_RDD0
                      : SINTCCMAPR10NoCE0ARA0RRh10hold): 1'bx))))) && !xpc10_stall)  TClo6_9_V_2 <= ((A_sA_SINT_CC_SCALbx22_ARB0[TClo6_9_V_0
                          ]==2'd3/*MS*/)? ((xpc10nz==8'd237/*US*/)? A_SINT_CC_MAPR12NoCE3_ARB0_RDD0: SINTCCMAPR12NoCE3ARB0RRh10hold): ((A_sA_SINT_CC_SCALbx22_ARB0
                          [TClo6_9_V_0]==2'd2/*MS*/)? ((xpc10nz==8'd237/*US*/)? A_SINT_CC_MAPR12NoCE2_ARB0_RDD0: SINTCCMAPR12NoCE2ARB0RRh10hold
                          ): ((A_sA_SINT_CC_SCALbx22_ARB0[TClo6_9_V_0]==1'd1/*MS*/)? ((xpc10nz==8'd237/*US*/)? A_SINT_CC_MAPR12NoCE1_ARB0_RDD0
                          : SINTCCMAPR12NoCE1ARB0RRh10hold): ((A_sA_SINT_CC_SCALbx22_ARB0[TClo6_9_V_0]==0/*MS*/)? ((xpc10nz==8'd237/*US*/)? A_SINT_CC_MAPR12NoCE0_ARB0_RDD0
                          : SINTCCMAPR12NoCE0ARB0RRh10hold): 32'bx))));

                          if ((TTMT4Main_V_11!=((A_sA_SINT_CC_SCALbx20_ARA0[TClo6_9_V_0]==2'd3/*MS*/)? ((xpc10nz==8'd237/*US*/)? A_SINT_CC_MAPR10NoCE3_ARA0_RDD0
                      : SINTCCMAPR10NoCE3ARA0RRh10hold): ((A_sA_SINT_CC_SCALbx20_ARA0[TClo6_9_V_0]==2'd2/*MS*/)? ((xpc10nz==8'd237/*US*/)? A_SINT_CC_MAPR10NoCE2_ARA0_RDD0
                      : SINTCCMAPR10NoCE2ARA0RRh10hold): ((A_sA_SINT_CC_SCALbx20_ARA0[TClo6_9_V_0]==1'd1/*MS*/)? ((xpc10nz==8'd237/*US*/)? A_SINT_CC_MAPR10NoCE1_ARA0_RDD0
                      : SINTCCMAPR10NoCE1ARA0RRh10hold): ((A_sA_SINT_CC_SCALbx20_ARA0[TClo6_9_V_0]==0/*MS*/)? ((xpc10nz==8'd237/*US*/)? A_SINT_CC_MAPR10NoCE0_ARA0_RDD0
                      : SINTCCMAPR10NoCE0ARA0RRh10hold): 1'bx))))) && !xpc10_stall)  TClo6_9_V_0 <= 32'd1+TClo6_9_V_0;
                          if ((TClo6_9_V_0==3'd4/*US*/) && (TTMT4Main_V_11==((A_sA_SINT_CC_SCALbx20_ARA0[TClo6_9_V_0]==2'd3/*MS*/)? ((xpc10nz
                      ==8'd237/*US*/)? A_SINT_CC_MAPR10NoCE3_ARA0_RDD0: SINTCCMAPR10NoCE3ARA0RRh10hold): ((A_sA_SINT_CC_SCALbx20_ARA0
                      [TClo6_9_V_0]==2'd2/*MS*/)? ((xpc10nz==8'd237/*US*/)? A_SINT_CC_MAPR10NoCE2_ARA0_RDD0: SINTCCMAPR10NoCE2ARA0RRh10hold
                      ): ((A_sA_SINT_CC_SCALbx20_ARA0[TClo6_9_V_0]==1'd1/*MS*/)? ((xpc10nz==8'd237/*US*/)? A_SINT_CC_MAPR10NoCE1_ARA0_RDD0
                      : SINTCCMAPR10NoCE1ARA0RRh10hold): ((A_sA_SINT_CC_SCALbx20_ARA0[TClo6_9_V_0]==0/*MS*/)? ((xpc10nz==8'd237/*US*/)? A_SINT_CC_MAPR10NoCE0_ARA0_RDD0
                      : SINTCCMAPR10NoCE0ARA0RRh10hold): 1'bx))))))  xpc10nz <= 8'd238/*xpc10nz*/;
                          if ((TClo6_9_V_0!=3'd4/*US*/) && (TTMT4Main_V_11==((A_sA_SINT_CC_SCALbx20_ARA0[TClo6_9_V_0]==2'd3/*MS*/)? ((xpc10nz
                      ==8'd237/*US*/)? A_SINT_CC_MAPR10NoCE3_ARA0_RDD0: SINTCCMAPR10NoCE3ARA0RRh10hold): ((A_sA_SINT_CC_SCALbx20_ARA0
                      [TClo6_9_V_0]==2'd2/*MS*/)? ((xpc10nz==8'd237/*US*/)? A_SINT_CC_MAPR10NoCE2_ARA0_RDD0: SINTCCMAPR10NoCE2ARA0RRh10hold
                      ): ((A_sA_SINT_CC_SCALbx20_ARA0[TClo6_9_V_0]==1'd1/*MS*/)? ((xpc10nz==8'd237/*US*/)? A_SINT_CC_MAPR10NoCE1_ARA0_RDD0
                      : SINTCCMAPR10NoCE1ARA0RRh10hold): ((A_sA_SINT_CC_SCALbx20_ARA0[TClo6_9_V_0]==0/*MS*/)? ((xpc10nz==8'd237/*US*/)? A_SINT_CC_MAPR10NoCE0_ARA0_RDD0
                      : SINTCCMAPR10NoCE0ARA0RRh10hold): 1'bx))))))  xpc10nz <= 8'd239/*xpc10nz*/;
                          if ((TTMT4Main_V_11!=((A_sA_SINT_CC_SCALbx20_ARA0[TClo6_9_V_0]==2'd3/*MS*/)? ((xpc10nz==8'd237/*US*/)? A_SINT_CC_MAPR10NoCE3_ARA0_RDD0
                      : SINTCCMAPR10NoCE3ARA0RRh10hold): ((A_sA_SINT_CC_SCALbx20_ARA0[TClo6_9_V_0]==2'd2/*MS*/)? ((xpc10nz==8'd237/*US*/)? A_SINT_CC_MAPR10NoCE2_ARA0_RDD0
                      : SINTCCMAPR10NoCE2ARA0RRh10hold): ((A_sA_SINT_CC_SCALbx20_ARA0[TClo6_9_V_0]==1'd1/*MS*/)? ((xpc10nz==8'd237/*US*/)? A_SINT_CC_MAPR10NoCE1_ARA0_RDD0
                      : SINTCCMAPR10NoCE1ARA0RRh10hold): ((A_sA_SINT_CC_SCALbx20_ARA0[TClo6_9_V_0]==0/*MS*/)? ((xpc10nz==8'd237/*US*/)? A_SINT_CC_MAPR10NoCE0_ARA0_RDD0
                      : SINTCCMAPR10NoCE0ARA0RRh10hold): 1'bx))))))  xpc10nz <= 8'd242/*xpc10nz*/;
                           end 
                      
                  8'd242/*US*/:  begin 
                      if ((TClo6_9_V_0<3'd4) && (TClo6_9_V_0==3'd4/*US*/))  begin 
                               A_SINT_CC_SCALbx24_stats_lookup_probes <= 32'd1+A_SINT_CC_SCALbx24_stats_lookup_probes;
                               TTMT4Main_V_14 <= -32'h5;
                               TCl6_SPILL_256 <= -32'd5;
                               end 
                              if ((TClo6_9_V_0==3'd4/*US*/) && !xpc10_stall)  begin 
                               TTMT4Main_V_14 <= -32'h5;
                               TCl6_SPILL_256 <= -32'd5;
                               end 
                              if ((TClo6_9_V_0<3'd4) && !xpc10_stall)  A_SINT_CC_SCALbx24_stats_lookup_probes <= 32'd1+A_SINT_CC_SCALbx24_stats_lookup_probes
                          ;

                          if ((TClo6_9_V_0==3'd4/*US*/))  xpc10nz <= 8'd238/*xpc10nz*/;
                          if ((TClo6_9_V_0>=3'd4) && (TClo6_9_V_0!=3'd4/*US*/))  xpc10nz <= 8'd243/*xpc10nz*/;
                          if ((TClo6_9_V_0<3'd4))  xpc10nz <= 7'd105/*xpc10nz*/;
                           end 
                      
                  8'd249/*US*/:  begin 
                      if (!(!TCin1_9_V_0) && (A_SINT_CC_SCALbx24_next_free==3'd4*A_SINT_CC_SCALbx24_waycap) && !xpc10_stall)  begin 
                               TCi1_SPILL_256 <= -32'd2;
                               TTMT4Main_V_7 <= -32'h2;
                               end 
                              if (!TCin1_9_V_0 && !xpc10_stall)  begin 
                               TCi1_SPILL_256 <= -32'd4;
                               TTMT4Main_V_7 <= -32'h4;
                               end 
                              if (!(!TCin1_9_V_0) && (A_SINT_CC_SCALbx24_next_free!=3'd4*A_SINT_CC_SCALbx24_waycap) && !xpc10_stall) 
                       fastspilldup16 <= A_SINT_CC_SCALbx24_next_free;
                          if ((!(!TCin1_9_V_0)? (A_SINT_CC_SCALbx24_next_free==3'd4*A_SINT_CC_SCALbx24_waycap): 1'd1))  xpc10nz <= 8'd250
                          /*xpc10nz*/;

                          if (!(!TCin1_9_V_0) && (A_SINT_CC_SCALbx24_next_free!=3'd4*A_SINT_CC_SCALbx24_waycap))  xpc10nz <= 8'd254/*xpc10nz*/;
                           end 
                      
                  9'd259/*US*/:  begin 
                      if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=1'd1/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=1'd1/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=0/*MS*/) && !xpc10_stall)  begin 
                               TCi1_SPILL_256 <= 32'd0;
                               TTMT4Main_V_7 <= 32'h0;
                               end 
                              if ((TCin1_9_V_4<3'd4) && (TCin1_9_V_4==3'd4/*US*/))  begin 
                               A_SINT_CC_SCALbx24_stats_insert_probes <= 32'd1+A_SINT_CC_SCALbx24_stats_insert_probes;
                               TCin1_9_V_1 <= 32'd1+TCin1_9_V_1;
                               end 
                              if ((TCin1_9_V_4<3'd4))  xpc10nz <= 9'd341/*xpc10nz*/;
                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=1'd1/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=1'd1/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=0/*MS*/))  xpc10nz <= 8'd250/*xpc10nz*/;
                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=1'd1/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==0/*MS*/))  xpc10nz
                           <= 9'd283/*xpc10nz*/;

                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=1'd1/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==1'd1/*MS*/))  xpc10nz
                           <= 9'd282/*xpc10nz*/;

                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=1'd1/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd2/*MS*/))  xpc10nz
                           <= 9'd281/*xpc10nz*/;

                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=1'd1/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd3/*MS*/))  xpc10nz
                           <= 9'd280/*xpc10nz*/;

                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==0/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd2/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=0/*MS*/))  xpc10nz
                           <= 9'd279/*xpc10nz*/;

                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==0/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==0/*MS*/))  xpc10nz <= 9'd278/*xpc10nz*/;
                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==0/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==1'd1/*MS*/))  xpc10nz <= 9'd277/*xpc10nz*/;
                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==0/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd2/*MS*/))  xpc10nz <= 9'd276/*xpc10nz*/;
                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==0/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd3/*MS*/))  xpc10nz <= 9'd275/*xpc10nz*/;
                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==1'd1/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd2/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=0/*MS*/))  xpc10nz
                           <= 9'd274/*xpc10nz*/;

                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==1'd1/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==0/*MS*/))  xpc10nz <= 9'd273/*xpc10nz*/;
                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==1'd1/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==1'd1/*MS*/))  xpc10nz <= 9'd272/*xpc10nz*/;
                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==1'd1/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd2/*MS*/))  xpc10nz <= 9'd271/*xpc10nz*/;
                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==1'd1/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd3/*MS*/))  xpc10nz <= 9'd270/*xpc10nz*/;
                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd2/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd2/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=0/*MS*/))  xpc10nz
                           <= 9'd269/*xpc10nz*/;

                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd2/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==0/*MS*/))  xpc10nz <= 9'd268/*xpc10nz*/;
                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd2/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==1'd1/*MS*/))  xpc10nz <= 9'd267/*xpc10nz*/;
                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd2/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd2/*MS*/))  xpc10nz <= 9'd266/*xpc10nz*/;
                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd2/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd3/*MS*/))  xpc10nz <= 9'd265/*xpc10nz*/;
                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd2/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=0/*MS*/))  xpc10nz
                           <= 9'd264/*xpc10nz*/;

                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==0/*MS*/))  xpc10nz <= 9'd263/*xpc10nz*/;
                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==1'd1/*MS*/))  xpc10nz <= 9'd262/*xpc10nz*/;
                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd2/*MS*/))  xpc10nz <= 9'd261/*xpc10nz*/;
                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd3/*MS*/))  xpc10nz <= 9'd260/*xpc10nz*/;
                          if ((TCin1_9_V_4==3'd4/*US*/))  xpc10nz <= 9'd284/*xpc10nz*/;
                          if ((TCin1_9_V_4<3'd4) && !xpc10_stall)  A_SINT_CC_SCALbx24_stats_insert_probes <= 32'd1+A_SINT_CC_SCALbx24_stats_insert_probes
                          ;

                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=1'd1/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==0/*MS*/) && !xpc10_stall
                      )  TCi1_SPILL_256 <= 32'd0;
                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=1'd1/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==1'd1/*MS*/) && 
                      !xpc10_stall)  TCi1_SPILL_256 <= 32'd0;
                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=1'd1/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd2/*MS*/) && 
                      !xpc10_stall)  TCi1_SPILL_256 <= 32'd0;
                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=1'd1/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd3/*MS*/) && 
                      !xpc10_stall)  TCi1_SPILL_256 <= 32'd0;
                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==0/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd2/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=0/*MS*/) && 
                      !xpc10_stall)  TCi1_SPILL_256 <= 32'd0;
                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==1'd1/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd2/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=0/*MS*/) && 
                      !xpc10_stall)  TCi1_SPILL_256 <= 32'd0;
                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd2/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd2/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=0/*MS*/) && 
                      !xpc10_stall)  TCi1_SPILL_256 <= 32'd0;
                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd2/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=0/*MS*/) && 
                      !xpc10_stall)  TCi1_SPILL_256 <= 32'd0;
                          if ((TCin1_9_V_4==3'd4/*US*/) && !xpc10_stall)  TCin1_9_V_1 <= 32'd1+TCin1_9_V_1;
                           end 
                      
                  9'd289/*US*/:  begin 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim
                      ]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [A_SINT_CC_SCALbx24_next_victim]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]!=2'd3
                      /*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [A_SINT_CC_SCALbx24_next_victim]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]!=0
                      /*MS*/) && !xpc10_stall)  begin 
                               TCin1_9_V_2 <= TCin1_9_V_7;
                               TCin1_9_V_0 <= TCin1_9_V_6;
                               end 
                              if ((A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]==2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [A_SINT_CC_SCALbx24_next_victim]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]!=2'd2
                      /*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [A_SINT_CC_SCALbx24_next_victim]!=0/*MS*/) && !xpc10_stall)  TCin1_9_V_0 <= TCin1_9_V_6;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]==2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [A_SINT_CC_SCALbx24_next_victim]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]!=2'd2
                      /*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [A_SINT_CC_SCALbx24_next_victim]!=0/*MS*/) && !xpc10_stall)  TCin1_9_V_0 <= TCin1_9_V_6;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]==1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [A_SINT_CC_SCALbx24_next_victim]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]!=2'd2
                      /*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [A_SINT_CC_SCALbx24_next_victim]!=0/*MS*/) && !xpc10_stall)  TCin1_9_V_0 <= TCin1_9_V_6;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]==0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim
                      ]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [A_SINT_CC_SCALbx24_next_victim]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]!=0
                      /*MS*/) && !xpc10_stall)  TCin1_9_V_0 <= TCin1_9_V_6;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [A_SINT_CC_SCALbx24_next_victim]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]!=1'd1
                      /*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [A_SINT_CC_SCALbx24_next_victim]==2'd3/*MS*/) && !xpc10_stall)  TCin1_9_V_0 <= TCin1_9_V_6;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [A_SINT_CC_SCALbx24_next_victim]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]!=1'd1
                      /*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [A_SINT_CC_SCALbx24_next_victim]==2'd2/*MS*/) && !xpc10_stall)  TCin1_9_V_0 <= TCin1_9_V_6;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [A_SINT_CC_SCALbx24_next_victim]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]!=1'd1
                      /*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [A_SINT_CC_SCALbx24_next_victim]==1'd1/*MS*/) && !xpc10_stall)  TCin1_9_V_0 <= TCin1_9_V_6;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [A_SINT_CC_SCALbx24_next_victim]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]!=1'd1
                      /*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [A_SINT_CC_SCALbx24_next_victim]==0/*MS*/) && !xpc10_stall)  TCin1_9_V_0 <= TCin1_9_V_6;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]==2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [A_SINT_CC_SCALbx24_next_victim]==2'd3/*MS*/))  xpc10nz <= 9'd290/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]==2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [A_SINT_CC_SCALbx24_next_victim]==2'd2/*MS*/))  xpc10nz <= 9'd291/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]==2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [A_SINT_CC_SCALbx24_next_victim]==1'd1/*MS*/))  xpc10nz <= 9'd292/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]==2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [A_SINT_CC_SCALbx24_next_victim]==0/*MS*/))  xpc10nz <= 9'd293/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]==2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [A_SINT_CC_SCALbx24_next_victim]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]!=2'd2
                      /*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [A_SINT_CC_SCALbx24_next_victim]!=0/*MS*/))  xpc10nz <= 9'd294/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]==2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [A_SINT_CC_SCALbx24_next_victim]==2'd3/*MS*/))  xpc10nz <= 9'd295/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]==2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [A_SINT_CC_SCALbx24_next_victim]==2'd2/*MS*/))  xpc10nz <= 9'd296/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]==2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [A_SINT_CC_SCALbx24_next_victim]==1'd1/*MS*/))  xpc10nz <= 9'd297/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]==2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [A_SINT_CC_SCALbx24_next_victim]==0/*MS*/))  xpc10nz <= 9'd298/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]==2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [A_SINT_CC_SCALbx24_next_victim]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]!=2'd2
                      /*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [A_SINT_CC_SCALbx24_next_victim]!=0/*MS*/))  xpc10nz <= 9'd299/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]==1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [A_SINT_CC_SCALbx24_next_victim]==2'd3/*MS*/))  xpc10nz <= 9'd300/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]==1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [A_SINT_CC_SCALbx24_next_victim]==2'd2/*MS*/))  xpc10nz <= 9'd301/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]==1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [A_SINT_CC_SCALbx24_next_victim]==1'd1/*MS*/))  xpc10nz <= 9'd302/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]==1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [A_SINT_CC_SCALbx24_next_victim]==0/*MS*/))  xpc10nz <= 9'd303/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]==1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [A_SINT_CC_SCALbx24_next_victim]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]!=2'd2
                      /*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [A_SINT_CC_SCALbx24_next_victim]!=0/*MS*/))  xpc10nz <= 9'd304/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]==0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim
                      ]==2'd3/*MS*/))  xpc10nz <= 9'd305/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]==0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim
                      ]==2'd2/*MS*/))  xpc10nz <= 9'd306/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]==0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim
                      ]==1'd1/*MS*/))  xpc10nz <= 9'd307/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]==0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim
                      ]==0/*MS*/))  xpc10nz <= 9'd308/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]==0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim
                      ]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [A_SINT_CC_SCALbx24_next_victim]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]!=0
                      /*MS*/))  xpc10nz <= 9'd309/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [A_SINT_CC_SCALbx24_next_victim]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]!=1'd1
                      /*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [A_SINT_CC_SCALbx24_next_victim]==2'd3/*MS*/))  xpc10nz <= 9'd310/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [A_SINT_CC_SCALbx24_next_victim]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]!=1'd1
                      /*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [A_SINT_CC_SCALbx24_next_victim]==2'd2/*MS*/))  xpc10nz <= 9'd311/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [A_SINT_CC_SCALbx24_next_victim]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]!=1'd1
                      /*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [A_SINT_CC_SCALbx24_next_victim]==1'd1/*MS*/))  xpc10nz <= 9'd312/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [A_SINT_CC_SCALbx24_next_victim]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]!=1'd1
                      /*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [A_SINT_CC_SCALbx24_next_victim]==0/*MS*/))  xpc10nz <= 9'd313/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [A_SINT_CC_SCALbx24_next_victim]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]!=1'd1
                      /*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[A_SINT_CC_SCALbx24_next_victim]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [A_SINT_CC_SCALbx24_next_victim]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]!=2'd2
                      /*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [A_SINT_CC_SCALbx24_next_victim]!=0/*MS*/))  xpc10nz <= 9'd323/*xpc10nz*/;
                           end 
                      
                  9'd314/*US*/:  begin 
                      if ((A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]==0/*MS*/))  xpc10nz <= 9'd317/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]==0/*MS*/) && !xpc10_stall)  TCin1_9_V_0 <= TCin1_9_V_6
                          ;

                          if ((A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]==1'd1/*MS*/))  xpc10nz <= 9'd316/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [A_SINT_CC_SCALbx24_next_victim]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]!=0
                      /*MS*/) && !xpc10_stall)  begin 
                               TCin1_9_V_2 <= TCin1_9_V_7;
                               TCin1_9_V_0 <= TCin1_9_V_6;
                               end 
                              if ((A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]==1'd1/*MS*/) && !xpc10_stall)  TCin1_9_V_0
                           <= TCin1_9_V_6;

                          if ((A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]==2'd2/*MS*/) && !xpc10_stall)  TCin1_9_V_0 <= TCin1_9_V_6
                          ;

                          if ((A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]==2'd2/*MS*/))  xpc10nz <= 9'd315/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [A_SINT_CC_SCALbx24_next_victim]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]!=0
                      /*MS*/))  xpc10nz <= 9'd323/*xpc10nz*/;
                           end 
                      
                  9'd324/*US*/:  begin 
                      if ((A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]==0/*MS*/))  xpc10nz <= 9'd326/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]==0/*MS*/) && !xpc10_stall)  TCin1_9_V_0 <= TCin1_9_V_6
                          ;

                          if ((A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]==1'd1/*MS*/))  xpc10nz <= 9'd325/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [A_SINT_CC_SCALbx24_next_victim]!=0/*MS*/) && !xpc10_stall)  begin 
                               TCin1_9_V_2 <= TCin1_9_V_7;
                               TCin1_9_V_0 <= TCin1_9_V_6;
                               end 
                              if ((A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]==1'd1/*MS*/) && !xpc10_stall)  TCin1_9_V_0
                           <= TCin1_9_V_6;

                          if ((A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [A_SINT_CC_SCALbx24_next_victim]!=0/*MS*/))  xpc10nz <= 9'd323/*xpc10nz*/;
                           end 
                      
                  9'd330/*US*/:  begin 
                      if ((A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==0/*MS*/))  xpc10nz <= 9'd333/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==0/*MS*/) && !xpc10_stall)  TCi1_SPILL_256 <= 32'd0;
                          if ((A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==1'd1/*MS*/))  xpc10nz <= 9'd332/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=1'd1
                      /*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=0/*MS*/) && !xpc10_stall)  begin 
                               TCi1_SPILL_256 <= 32'd0;
                               TTMT4Main_V_7 <= 32'h0;
                               end 
                              if ((A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==1'd1/*MS*/) && !xpc10_stall)  TCi1_SPILL_256 <= 32'd0;
                          if ((A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd2/*MS*/) && !xpc10_stall)  TCi1_SPILL_256 <= 32'd0;
                          if ((A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd2/*MS*/))  xpc10nz <= 9'd331/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=1'd1
                      /*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=0/*MS*/))  xpc10nz <= 8'd250/*xpc10nz*/;
                           end 
                      
                  9'd335/*US*/:  begin 
                      if ((A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==0/*MS*/))  xpc10nz <= 9'd337/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==0/*MS*/) && !xpc10_stall)  TCi1_SPILL_256 <= 32'd0;
                          if ((A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==1'd1/*MS*/))  xpc10nz <= 9'd336/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=0/*MS*/) && 
                      !xpc10_stall)  begin 
                               TCi1_SPILL_256 <= 32'd0;
                               TTMT4Main_V_7 <= 32'h0;
                               end 
                              if ((A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==1'd1/*MS*/) && !xpc10_stall)  TCi1_SPILL_256 <= 32'd0;
                          if ((A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=0/*MS*/)) 
                       xpc10nz <= 8'd250/*xpc10nz*/;
                           end 
                      
                  9'd473/*US*/:  begin 
                      if ((TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [TCin1_9_V_4]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [TCin1_9_V_4]!=0/*MS*/) && !xpc10_stall)  begin 
                               TCi1_SPILL_256 <= 32'd0;
                               TTMT4Main_V_7 <= 32'h0;
                               end 
                              if ((TCin1_9_V_4==3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [TCin1_9_V_4]!=0/*MS*/) && !xpc10_stall)  TCin1_9_V_1 <= 32'd1+TCin1_9_V_1;
                          if (((xpc10nz==9'd473/*US*/)? !A_SINT_CC_MAPR10NoCE3_ARA0_RDD0 && !xpc10_stall: !SINTCCMAPR10NoCE3ARA0RRh10hold
                       && !xpc10_stall) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4
                      ]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4
                      ]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd3/*MS*/) && (TCin1_9_V_4!=3'd4/*US*/))  TCi1_SPILL_256
                           <= 32'd0;

                          if (((xpc10nz==9'd473/*US*/)? !A_SINT_CC_MAPR10NoCE2_ARA0_RDD0 && !xpc10_stall: !SINTCCMAPR10NoCE2ARA0RRh10hold
                       && !xpc10_stall) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4
                      ]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4
                      ]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd2/*MS*/) && (TCin1_9_V_4!=3'd4/*US*/))  TCi1_SPILL_256
                           <= 32'd0;

                          if (((xpc10nz==9'd473/*US*/)? !A_SINT_CC_MAPR10NoCE1_ARA0_RDD0 && !xpc10_stall: !SINTCCMAPR10NoCE1ARA0RRh10hold
                       && !xpc10_stall) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4
                      ]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4
                      ]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==1'd1/*MS*/) && (TCin1_9_V_4!=3'd4/*US*/))  TCi1_SPILL_256
                           <= 32'd0;

                          if (((xpc10nz==9'd473/*US*/)? !A_SINT_CC_MAPR10NoCE0_ARA0_RDD0 && !xpc10_stall: !SINTCCMAPR10NoCE0ARA0RRh10hold
                       && !xpc10_stall) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4
                      ]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4
                      ]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==0/*MS*/) && (TCin1_9_V_4!=3'd4/*US*/))  TCi1_SPILL_256
                           <= 32'd0;

                          if ((TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [TCin1_9_V_4]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd3/*MS*/) && !xpc10_stall)  TCi1_SPILL_256
                           <= 32'd0;

                          if ((TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [TCin1_9_V_4]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd2/*MS*/) && !xpc10_stall)  TCi1_SPILL_256
                           <= 32'd0;

                          if ((TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [TCin1_9_V_4]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==1'd1/*MS*/) && !xpc10_stall)  TCi1_SPILL_256
                           <= 32'd0;

                          if ((TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [TCin1_9_V_4]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==0/*MS*/) && !xpc10_stall)  TCi1_SPILL_256 <= 32'd0
                          ;

                          if (((xpc10nz==9'd473/*US*/)? (!(!A_SINT_CC_MAPR10NoCE0_ARA0_RDD0) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4
                      ]==0/*MS*/) || !(!A_SINT_CC_MAPR10NoCE1_ARA0_RDD0) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==1'd1/*MS*/) || 
                      !(!A_SINT_CC_MAPR10NoCE2_ARA0_RDD0) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd2/*MS*/) || !(!A_SINT_CC_MAPR10NoCE3_ARA0_RDD0
                      ) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd3/*MS*/)) && !xpc10_stall: (!(!SINTCCMAPR10NoCE0ARA0RRh10hold
                      ) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==0/*MS*/) || !(!SINTCCMAPR10NoCE1ARA0RRh10hold) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [TCin1_9_V_4]==1'd1/*MS*/) || !(!SINTCCMAPR10NoCE2ARA0RRh10hold) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd2
                      /*MS*/) || !(!SINTCCMAPR10NoCE3ARA0RRh10hold) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd3/*MS*/)) && !xpc10_stall
                      ))  TCin1_9_V_4 <= 32'd1+TCin1_9_V_4;
                          if (((xpc10nz==9'd473/*US*/)? !A_SINT_CC_MAPR10NoCE3_ARA0_RDD0: !SINTCCMAPR10NoCE3ARA0RRh10hold) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [TCin1_9_V_4]==2'd3/*MS*/) && (TCin1_9_V_4==3'd4/*US*/))  xpc10nz <= 9'd474/*xpc10nz*/;
                          if (((xpc10nz==9'd473/*US*/)? !A_SINT_CC_MAPR10NoCE3_ARA0_RDD0: !SINTCCMAPR10NoCE3ARA0RRh10hold) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [TCin1_9_V_4]==2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd3/*MS*/) && (TCin1_9_V_4!=3'd4/*US*/)) 
                       xpc10nz <= 9'd475/*xpc10nz*/;
                          if (((xpc10nz==9'd473/*US*/)? !A_SINT_CC_MAPR10NoCE3_ARA0_RDD0: !SINTCCMAPR10NoCE3ARA0RRh10hold) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [TCin1_9_V_4]==2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd3/*MS*/) && (TCin1_9_V_4!=3'd4/*US*/)) 
                       xpc10nz <= 9'd476/*xpc10nz*/;
                          if (((xpc10nz==9'd473/*US*/)? !A_SINT_CC_MAPR10NoCE3_ARA0_RDD0: !SINTCCMAPR10NoCE3ARA0RRh10hold) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [TCin1_9_V_4]==1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd3/*MS*/) && (TCin1_9_V_4!=3'd4/*US*/)) 
                       xpc10nz <= 9'd477/*xpc10nz*/;
                          if (((xpc10nz==9'd473/*US*/)? !A_SINT_CC_MAPR10NoCE3_ARA0_RDD0: !SINTCCMAPR10NoCE3ARA0RRh10hold) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [TCin1_9_V_4]==0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd3/*MS*/) && (TCin1_9_V_4!=3'd4/*US*/)) 
                       xpc10nz <= 9'd478/*xpc10nz*/;
                          if (((xpc10nz==9'd473/*US*/)? !A_SINT_CC_MAPR10NoCE3_ARA0_RDD0: !SINTCCMAPR10NoCE3ARA0RRh10hold) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [TCin1_9_V_4]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [TCin1_9_V_4]==2'd3/*MS*/) && (TCin1_9_V_4!=3'd4/*US*/))  xpc10nz <= 9'd479/*xpc10nz*/;
                          if (((xpc10nz==9'd473/*US*/)? !A_SINT_CC_MAPR10NoCE2_ARA0_RDD0: !SINTCCMAPR10NoCE2ARA0RRh10hold) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [TCin1_9_V_4]==2'd2/*MS*/) && (TCin1_9_V_4==3'd4/*US*/))  xpc10nz <= 9'd480/*xpc10nz*/;
                          if (((xpc10nz==9'd473/*US*/)? !A_SINT_CC_MAPR10NoCE2_ARA0_RDD0: !SINTCCMAPR10NoCE2ARA0RRh10hold) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [TCin1_9_V_4]==2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd2/*MS*/) && (TCin1_9_V_4!=3'd4/*US*/)) 
                       xpc10nz <= 9'd481/*xpc10nz*/;
                          if (((xpc10nz==9'd473/*US*/)? !A_SINT_CC_MAPR10NoCE2_ARA0_RDD0: !SINTCCMAPR10NoCE2ARA0RRh10hold) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [TCin1_9_V_4]==2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd2/*MS*/) && (TCin1_9_V_4!=3'd4/*US*/)) 
                       xpc10nz <= 9'd482/*xpc10nz*/;
                          if (((xpc10nz==9'd473/*US*/)? !A_SINT_CC_MAPR10NoCE2_ARA0_RDD0: !SINTCCMAPR10NoCE2ARA0RRh10hold) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [TCin1_9_V_4]==1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd2/*MS*/) && (TCin1_9_V_4!=3'd4/*US*/)) 
                       xpc10nz <= 9'd483/*xpc10nz*/;
                          if (((xpc10nz==9'd473/*US*/)? !A_SINT_CC_MAPR10NoCE2_ARA0_RDD0: !SINTCCMAPR10NoCE2ARA0RRh10hold) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [TCin1_9_V_4]==0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd2/*MS*/) && (TCin1_9_V_4!=3'd4/*US*/)) 
                       xpc10nz <= 9'd484/*xpc10nz*/;
                          if (((xpc10nz==9'd473/*US*/)? !A_SINT_CC_MAPR10NoCE2_ARA0_RDD0: !SINTCCMAPR10NoCE2ARA0RRh10hold) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [TCin1_9_V_4]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [TCin1_9_V_4]==2'd2/*MS*/) && (TCin1_9_V_4!=3'd4/*US*/))  xpc10nz <= 9'd485/*xpc10nz*/;
                          if (((xpc10nz==9'd473/*US*/)? !A_SINT_CC_MAPR10NoCE1_ARA0_RDD0: !SINTCCMAPR10NoCE1ARA0RRh10hold) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [TCin1_9_V_4]==1'd1/*MS*/) && (TCin1_9_V_4==3'd4/*US*/))  xpc10nz <= 9'd486/*xpc10nz*/;
                          if (((xpc10nz==9'd473/*US*/)? !A_SINT_CC_MAPR10NoCE1_ARA0_RDD0: !SINTCCMAPR10NoCE1ARA0RRh10hold) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [TCin1_9_V_4]==2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==1'd1/*MS*/) && (TCin1_9_V_4!=3'd4/*US*/)) 
                       xpc10nz <= 9'd487/*xpc10nz*/;
                          if (((xpc10nz==9'd473/*US*/)? !A_SINT_CC_MAPR10NoCE1_ARA0_RDD0: !SINTCCMAPR10NoCE1ARA0RRh10hold) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [TCin1_9_V_4]==2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==1'd1/*MS*/) && (TCin1_9_V_4!=3'd4/*US*/)) 
                       xpc10nz <= 9'd488/*xpc10nz*/;
                          if (((xpc10nz==9'd473/*US*/)? !A_SINT_CC_MAPR10NoCE1_ARA0_RDD0: !SINTCCMAPR10NoCE1ARA0RRh10hold) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [TCin1_9_V_4]==1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==1'd1/*MS*/) && (TCin1_9_V_4!=3'd4/*US*/)) 
                       xpc10nz <= 9'd489/*xpc10nz*/;
                          if (((xpc10nz==9'd473/*US*/)? !A_SINT_CC_MAPR10NoCE1_ARA0_RDD0: !SINTCCMAPR10NoCE1ARA0RRh10hold) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [TCin1_9_V_4]==0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==1'd1/*MS*/) && (TCin1_9_V_4!=3'd4/*US*/)) 
                       xpc10nz <= 9'd490/*xpc10nz*/;
                          if (((xpc10nz==9'd473/*US*/)? !A_SINT_CC_MAPR10NoCE1_ARA0_RDD0: !SINTCCMAPR10NoCE1ARA0RRh10hold) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [TCin1_9_V_4]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [TCin1_9_V_4]==1'd1/*MS*/) && (TCin1_9_V_4!=3'd4/*US*/))  xpc10nz <= 9'd491/*xpc10nz*/;
                          if (((xpc10nz==9'd473/*US*/)? !A_SINT_CC_MAPR10NoCE0_ARA0_RDD0: !SINTCCMAPR10NoCE0ARA0RRh10hold) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [TCin1_9_V_4]==0/*MS*/) && (TCin1_9_V_4==3'd4/*US*/))  xpc10nz <= 9'd492/*xpc10nz*/;
                          if (((xpc10nz==9'd473/*US*/)? !A_SINT_CC_MAPR10NoCE0_ARA0_RDD0: !SINTCCMAPR10NoCE0ARA0RRh10hold) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [TCin1_9_V_4]==2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==0/*MS*/) && (TCin1_9_V_4!=3'd4/*US*/)) 
                       xpc10nz <= 9'd493/*xpc10nz*/;
                          if (((xpc10nz==9'd473/*US*/)? !A_SINT_CC_MAPR10NoCE0_ARA0_RDD0: !SINTCCMAPR10NoCE0ARA0RRh10hold) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [TCin1_9_V_4]==2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==0/*MS*/) && (TCin1_9_V_4!=3'd4/*US*/)) 
                       xpc10nz <= 9'd494/*xpc10nz*/;
                          if (((xpc10nz==9'd473/*US*/)? !A_SINT_CC_MAPR10NoCE0_ARA0_RDD0: !SINTCCMAPR10NoCE0ARA0RRh10hold) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [TCin1_9_V_4]==1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==0/*MS*/) && (TCin1_9_V_4!=3'd4/*US*/)) 
                       xpc10nz <= 9'd495/*xpc10nz*/;
                          if (((xpc10nz==9'd473/*US*/)? !A_SINT_CC_MAPR10NoCE0_ARA0_RDD0: !SINTCCMAPR10NoCE0ARA0RRh10hold) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [TCin1_9_V_4]==0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==0/*MS*/) && (TCin1_9_V_4!=3'd4/*US*/))  xpc10nz
                           <= 9'd496/*xpc10nz*/;

                          if (((xpc10nz==9'd473/*US*/)? !A_SINT_CC_MAPR10NoCE0_ARA0_RDD0: !SINTCCMAPR10NoCE0ARA0RRh10hold) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [TCin1_9_V_4]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [TCin1_9_V_4]==0/*MS*/) && (TCin1_9_V_4!=3'd4/*US*/))  xpc10nz <= 9'd497/*xpc10nz*/;
                          if ((TCin1_9_V_4==3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [TCin1_9_V_4]!=0/*MS*/))  xpc10nz <= 9'd284/*xpc10nz*/;
                          if ((TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [TCin1_9_V_4]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd3/*MS*/))  xpc10nz <= 9'd498/*xpc10nz*/;
                          if ((TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [TCin1_9_V_4]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd2/*MS*/))  xpc10nz <= 9'd499/*xpc10nz*/;
                          if ((TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [TCin1_9_V_4]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==1'd1/*MS*/))  xpc10nz <= 9'd500/*xpc10nz*/;
                          if ((TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [TCin1_9_V_4]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==0/*MS*/))  xpc10nz <= 9'd501/*xpc10nz*/;
                          if ((TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [TCin1_9_V_4]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0
                      [TCin1_9_V_4]!=0/*MS*/))  xpc10nz <= 8'd250/*xpc10nz*/;
                          if (((xpc10nz==9'd473/*US*/)? !(!A_SINT_CC_MAPR10NoCE0_ARA0_RDD0) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4
                      ]==0/*MS*/) || !(!A_SINT_CC_MAPR10NoCE1_ARA0_RDD0) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==1'd1/*MS*/) || 
                      !(!A_SINT_CC_MAPR10NoCE2_ARA0_RDD0) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd2/*MS*/) || !(!A_SINT_CC_MAPR10NoCE3_ARA0_RDD0
                      ) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd3/*MS*/): !(!SINTCCMAPR10NoCE0ARA0RRh10hold) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [TCin1_9_V_4]==0/*MS*/) || !(!SINTCCMAPR10NoCE1ARA0RRh10hold) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==1'd1
                      /*MS*/) || !(!SINTCCMAPR10NoCE2ARA0RRh10hold) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd2/*MS*/) || !(!SINTCCMAPR10NoCE3ARA0RRh10hold
                      ) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd3/*MS*/)))  xpc10nz <= 9'd503/*xpc10nz*/;
                           end 
                      
                  9'd503/*US*/:  begin 
                      if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=1'd1/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=1'd1/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=0/*MS*/) && !xpc10_stall)  begin 
                               TCi1_SPILL_256 <= 32'd0;
                               TTMT4Main_V_7 <= 32'h0;
                               end 
                              if ((TCin1_9_V_4<3'd4) && (TCin1_9_V_4==3'd4/*US*/))  begin 
                               A_SINT_CC_SCALbx24_stats_insert_probes <= 32'd1+A_SINT_CC_SCALbx24_stats_insert_probes;
                               TCin1_9_V_1 <= 32'd1+TCin1_9_V_1;
                               end 
                              if ((TCin1_9_V_4<3'd4))  xpc10nz <= 9'd341/*xpc10nz*/;
                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=1'd1/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=1'd1/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=0/*MS*/))  xpc10nz <= 8'd250/*xpc10nz*/;
                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=1'd1/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==0/*MS*/))  xpc10nz
                           <= 10'd527/*xpc10nz*/;

                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=1'd1/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==1'd1/*MS*/))  xpc10nz
                           <= 10'd526/*xpc10nz*/;

                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=1'd1/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd2/*MS*/))  xpc10nz
                           <= 10'd525/*xpc10nz*/;

                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=1'd1/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd3/*MS*/))  xpc10nz
                           <= 10'd524/*xpc10nz*/;

                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==0/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd2/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=0/*MS*/))  xpc10nz
                           <= 10'd523/*xpc10nz*/;

                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==0/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==0/*MS*/))  xpc10nz <= 10'd522/*xpc10nz*/;
                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==0/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==1'd1/*MS*/))  xpc10nz <= 10'd521/*xpc10nz*/;
                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==0/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd2/*MS*/))  xpc10nz <= 10'd520/*xpc10nz*/;
                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==0/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd3/*MS*/))  xpc10nz <= 10'd519/*xpc10nz*/;
                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==1'd1/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd2/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=0/*MS*/))  xpc10nz
                           <= 10'd518/*xpc10nz*/;

                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==1'd1/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==0/*MS*/))  xpc10nz <= 10'd517/*xpc10nz*/;
                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==1'd1/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==1'd1/*MS*/))  xpc10nz <= 10'd516/*xpc10nz*/;
                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==1'd1/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd2/*MS*/))  xpc10nz <= 10'd515/*xpc10nz*/;
                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==1'd1/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd3/*MS*/))  xpc10nz <= 10'd514/*xpc10nz*/;
                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd2/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd2/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=0/*MS*/))  xpc10nz
                           <= 10'd513/*xpc10nz*/;

                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd2/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==0/*MS*/))  xpc10nz <= 10'd512/*xpc10nz*/;
                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd2/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==1'd1/*MS*/))  xpc10nz <= 9'd511/*xpc10nz*/;
                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd2/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd2/*MS*/))  xpc10nz <= 9'd510/*xpc10nz*/;
                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd2/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd3/*MS*/))  xpc10nz <= 9'd509/*xpc10nz*/;
                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd2/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=0/*MS*/))  xpc10nz
                           <= 9'd508/*xpc10nz*/;

                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==0/*MS*/))  xpc10nz <= 9'd507/*xpc10nz*/;
                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==1'd1/*MS*/))  xpc10nz <= 9'd506/*xpc10nz*/;
                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd2/*MS*/))  xpc10nz <= 9'd505/*xpc10nz*/;
                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd3/*MS*/))  xpc10nz <= 9'd504/*xpc10nz*/;
                          if ((TCin1_9_V_4==3'd4/*US*/))  xpc10nz <= 9'd284/*xpc10nz*/;
                          if ((TCin1_9_V_4<3'd4) && !xpc10_stall)  A_SINT_CC_SCALbx24_stats_insert_probes <= 32'd1+A_SINT_CC_SCALbx24_stats_insert_probes
                          ;

                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=1'd1/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==0/*MS*/) && !xpc10_stall
                      )  TCi1_SPILL_256 <= 32'd0;
                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=1'd1/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==1'd1/*MS*/) && 
                      !xpc10_stall)  TCi1_SPILL_256 <= 32'd0;
                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=1'd1/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd2/*MS*/) && 
                      !xpc10_stall)  TCi1_SPILL_256 <= 32'd0;
                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=1'd1/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==2'd3/*MS*/) && 
                      !xpc10_stall)  TCi1_SPILL_256 <= 32'd0;
                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==0/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd2/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=0/*MS*/) && 
                      !xpc10_stall)  TCi1_SPILL_256 <= 32'd0;
                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==1'd1/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd2/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=0/*MS*/) && 
                      !xpc10_stall)  TCi1_SPILL_256 <= 32'd0;
                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd2/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd2/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=0/*MS*/) && 
                      !xpc10_stall)  TCi1_SPILL_256 <= 32'd0;
                          if ((TCin1_9_V_4>=3'd4) && (TCin1_9_V_4!=3'd4/*US*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCin1_9_V_4]==2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=2'd2/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=0/*MS*/) && 
                      !xpc10_stall)  TCi1_SPILL_256 <= 32'd0;
                          if ((TCin1_9_V_4==3'd4/*US*/) && !xpc10_stall)  TCin1_9_V_1 <= 32'd1+TCin1_9_V_1;
                           end 
                      
                  10'd528/*US*/:  begin 
                      
                      case (A_sA_SINT_CC_SCALbx20_ARA0[TCCl0_12_V_1]) // synthesis full_case 
                          0/*MS*/:  xpc10nz <= 10'd531/*xpc10nz*/;

                          1'd1/*MS*/:  xpc10nz <= 10'd530/*xpc10nz*/;
                      endcase
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[TCCl0_12_V_1]==1'd1/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd1+TCCl0_12_V_1
                          ;

                          if ((A_sA_SINT_CC_SCALbx20_ARA0[TCCl0_12_V_1]==2'd2/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd1+TCCl0_12_V_1
                          ;

                          if (((A_sA_SINT_CC_SCALbx20_ARA0[TCCl0_12_V_1]==0/*MS*/)? !xpc10_stall: (A_sA_SINT_CC_SCALbx20_ARA0[TCCl0_12_V_1
                      ]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCCl0_12_V_1]!=1'd1/*MS*/) && !xpc10_stall))  TCCl0_12_V_1 <= 32'd1
                          +TCCl0_12_V_1;

                          if ((A_sA_SINT_CC_SCALbx20_ARA0[TCCl0_12_V_1]==2'd2/*MS*/))  xpc10nz <= 10'd529/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[TCCl0_12_V_1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCCl0_12_V_1]!=1'd1
                      /*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCCl0_12_V_1]!=0/*MS*/))  xpc10nz <= 10'd532/*xpc10nz*/;
                           end 
                      
                  10'd540/*US*/:  begin 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==0/*MS*/))  xpc10nz <= 10'd543/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==0/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd4;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==1'd1/*MS*/))  xpc10nz <= 10'd542/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==1'd1/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd4;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==2'd2/*MS*/))  xpc10nz <= 10'd541/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==2'd2/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd4;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd3]!=0/*MS*/) && !xpc10_stall)  begin 
                               TCCl0_12_V_0 <= 32'd1+TCCl0_12_V_0;
                               TCCl0_12_V_1 <= 32'd4;
                               end 
                              if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=1'd1/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=0/*MS*/))  xpc10nz <= 7'd65/*xpc10nz*/;
                           end 
                      
                  10'd544/*US*/:  begin 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==0/*MS*/))  xpc10nz <= 10'd546/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==0/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd4;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==1'd1/*MS*/))  xpc10nz <= 10'd545/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==1'd1/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd4;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=0/*MS*/) && !xpc10_stall
                      )  begin 
                               TCCl0_12_V_0 <= 32'd1+TCCl0_12_V_0;
                               TCCl0_12_V_1 <= 32'd4;
                               end 
                              if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=0/*MS*/))  xpc10nz
                           <= 7'd65/*xpc10nz*/;

                           end 
                      
                  10'd550/*US*/:  begin 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==0/*MS*/))  xpc10nz <= 10'd553/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==0/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd3;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==1'd1/*MS*/))  xpc10nz <= 10'd552/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==1'd1/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd3;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==2'd2/*MS*/))  xpc10nz <= 10'd551/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==2'd2/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd3;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=2'd2/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=0/*MS*/) && !xpc10_stall) 
                       begin 
                               TCCl0_12_V_0 <= 32'd1+TCCl0_12_V_0;
                               TCCl0_12_V_1 <= 32'd4;
                               end 
                              if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==2'd3/*MS*/) && !xpc10_stall) 
                       TCCl0_12_V_1 <= 32'd3;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==2'd2/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd3;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==1'd1/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd3;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==0/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd3;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==2'd3/*MS*/))  xpc10nz <= 10'd554/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==2'd2/*MS*/))  xpc10nz <= 10'd555/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==1'd1/*MS*/))  xpc10nz <= 10'd556/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==0/*MS*/))  xpc10nz <= 10'd557/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=2'd2/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=0/*MS*/))  xpc10nz <= 7'd65
                          /*xpc10nz*/;

                           end 
                      
                  10'd558/*US*/:  begin 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==0/*MS*/))  xpc10nz <= 10'd560/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==0/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd3;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==1'd1/*MS*/))  xpc10nz <= 10'd559/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==1'd1/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd3;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd3]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=1'd1
                      /*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=0/*MS*/) && !xpc10_stall)  begin 
                               TCCl0_12_V_0 <= 32'd1+TCCl0_12_V_0;
                               TCCl0_12_V_1 <= 32'd4;
                               end 
                              if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd3]==2'd3/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd3;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd3]==2'd2/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd3;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd3]==1'd1/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd3;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd3]==0/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd3;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd3]==2'd3/*MS*/))  xpc10nz <= 10'd561/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd3]==2'd2/*MS*/))  xpc10nz <= 10'd562/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd3]==1'd1/*MS*/))  xpc10nz <= 10'd563/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd3]==0/*MS*/))  xpc10nz <= 10'd564/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd3]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=1'd1
                      /*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=0/*MS*/))  xpc10nz <= 7'd65/*xpc10nz*/;
                           end 
                      
                  10'd565/*US*/:  begin 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==0/*MS*/))  xpc10nz <= 10'd566/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==0/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd3;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd3]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=0/*MS*/) && 
                      !xpc10_stall)  begin 
                               TCCl0_12_V_0 <= 32'd1+TCCl0_12_V_0;
                               TCCl0_12_V_1 <= 32'd4;
                               end 
                              if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==2'd3/*MS*/) && !xpc10_stall
                      )  TCCl0_12_V_1 <= 32'd3;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==2'd2/*MS*/) && !xpc10_stall
                      )  TCCl0_12_V_1 <= 32'd3;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==1'd1/*MS*/) && !xpc10_stall
                      )  TCCl0_12_V_1 <= 32'd3;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==0/*MS*/) && !xpc10_stall
                      )  TCCl0_12_V_1 <= 32'd3;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==2'd3/*MS*/))  xpc10nz
                           <= 10'd567/*xpc10nz*/;

                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==2'd2/*MS*/))  xpc10nz
                           <= 10'd568/*xpc10nz*/;

                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==1'd1/*MS*/))  xpc10nz
                           <= 10'd569/*xpc10nz*/;

                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==0/*MS*/))  xpc10nz <= 10'd570
                          /*xpc10nz*/;

                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd3]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=0/*MS*/)) 
                       xpc10nz <= 7'd65/*xpc10nz*/;
                           end 
                      
                  10'd571/*US*/:  begin 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==0/*MS*/))  xpc10nz <= 10'd575/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==0/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd3;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==1'd1/*MS*/))  xpc10nz <= 10'd574/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd3]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=0/*MS*/) && !xpc10_stall)  begin 
                               TCCl0_12_V_0 <= 32'd1+TCCl0_12_V_0;
                               TCCl0_12_V_1 <= 32'd4;
                               end 
                              if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==1'd1/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd3;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==2'd2/*MS*/))  xpc10nz <= 10'd573/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==2'd2/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd3;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd3]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=0/*MS*/))  xpc10nz <= 7'd65/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==2'd3/*MS*/))  xpc10nz <= 10'd572/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==2'd3/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd3;
                           end 
                      
                  10'd576/*US*/:  begin 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]==0/*MS*/))  xpc10nz <= 10'd579/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]==0/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd2;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]==1'd1/*MS*/))  xpc10nz <= 10'd578/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]==1'd1/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd2;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]==2'd2/*MS*/))  xpc10nz <= 10'd577/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd3]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=1'd1
                      /*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=0/*MS*/) && !xpc10_stall)  begin 
                               TCCl0_12_V_0 <= 32'd1+TCCl0_12_V_0;
                               TCCl0_12_V_1 <= 32'd4;
                               end 
                              if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]==2'd2/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd2;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==2'd3/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd2;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==2'd2/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd2;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==1'd1/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd2;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==0/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd2;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd3]==2'd3/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd3;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd3]==2'd2/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd3;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd3]==1'd1/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd3;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd3]==0/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd3;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==2'd3/*MS*/))  xpc10nz <= 10'd580/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==2'd2/*MS*/))  xpc10nz <= 10'd581/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==1'd1/*MS*/))  xpc10nz <= 10'd582/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==0/*MS*/))  xpc10nz <= 10'd583/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd3]==2'd3/*MS*/))  xpc10nz <= 10'd584/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd3]==2'd2/*MS*/))  xpc10nz <= 10'd585/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd3]==1'd1/*MS*/))  xpc10nz <= 10'd586/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd3]==0/*MS*/))  xpc10nz <= 10'd587/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd3]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=1'd1
                      /*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=0/*MS*/))  xpc10nz <= 7'd65/*xpc10nz*/;
                           end 
                      
                  10'd588/*US*/:  begin 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]==0/*MS*/))  xpc10nz <= 10'd590/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]==0/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd2;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]==1'd1/*MS*/))  xpc10nz <= 10'd589/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]==1'd1/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd2;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1
                      /*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd3]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=0/*MS*/) && 
                      !xpc10_stall)  begin 
                               TCCl0_12_V_0 <= 32'd1+TCCl0_12_V_0;
                               TCCl0_12_V_1 <= 32'd4;
                               end 
                              if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]==2'd3/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd2;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]==2'd2/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd2;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]==1'd1/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd2;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]==0/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd2;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1
                      /*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==2'd3/*MS*/) && !xpc10_stall
                      )  TCCl0_12_V_1 <= 32'd3;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1
                      /*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==2'd2/*MS*/) && !xpc10_stall
                      )  TCCl0_12_V_1 <= 32'd3;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1
                      /*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==1'd1/*MS*/) && !xpc10_stall
                      )  TCCl0_12_V_1 <= 32'd3;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1
                      /*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==0/*MS*/) && !xpc10_stall
                      )  TCCl0_12_V_1 <= 32'd3;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]==2'd3/*MS*/))  xpc10nz <= 10'd591/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]==2'd2/*MS*/))  xpc10nz <= 10'd592/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]==1'd1/*MS*/))  xpc10nz <= 10'd593/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]==0/*MS*/))  xpc10nz <= 10'd594/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1
                      /*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==2'd3/*MS*/))  xpc10nz
                           <= 10'd595/*xpc10nz*/;

                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1
                      /*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==2'd2/*MS*/))  xpc10nz
                           <= 10'd596/*xpc10nz*/;

                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1
                      /*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==1'd1/*MS*/))  xpc10nz
                           <= 10'd597/*xpc10nz*/;

                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1
                      /*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==0/*MS*/))  xpc10nz
                           <= 10'd598/*xpc10nz*/;

                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1
                      /*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd3]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=0/*MS*/)) 
                       xpc10nz <= 7'd65/*xpc10nz*/;
                           end 
                      
                  10'd599/*US*/:  begin 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]==0/*MS*/))  xpc10nz <= 10'd600/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]==0/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd2;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd3]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=0/*MS*/) && !xpc10_stall)  begin 
                               TCCl0_12_V_0 <= 32'd1+TCCl0_12_V_0;
                               TCCl0_12_V_1 <= 32'd4;
                               end 
                              if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==2'd3/*MS*/) && !xpc10_stall
                      )  TCCl0_12_V_1 <= 32'd2;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==2'd2/*MS*/) && !xpc10_stall
                      )  TCCl0_12_V_1 <= 32'd2;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==1'd1/*MS*/) && !xpc10_stall
                      )  TCCl0_12_V_1 <= 32'd2;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==0/*MS*/) && !xpc10_stall
                      )  TCCl0_12_V_1 <= 32'd2;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==2'd3/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd3;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==2'd2/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd3;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==1'd1/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd3;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==0/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd3;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==2'd3/*MS*/))  xpc10nz
                           <= 10'd601/*xpc10nz*/;

                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==2'd2/*MS*/))  xpc10nz
                           <= 10'd602/*xpc10nz*/;

                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==1'd1/*MS*/))  xpc10nz
                           <= 10'd603/*xpc10nz*/;

                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==0/*MS*/))  xpc10nz <= 10'd604
                          /*xpc10nz*/;

                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==2'd3/*MS*/))  xpc10nz <= 10'd605/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==2'd2/*MS*/))  xpc10nz <= 10'd606/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==1'd1/*MS*/))  xpc10nz <= 10'd607/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==0/*MS*/))  xpc10nz <= 10'd608/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[1'd1]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd3]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=0/*MS*/))  xpc10nz <= 7'd65/*xpc10nz*/;
                           end 
                      
                  10'd609/*US*/:  begin 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==0/*MS*/))  xpc10nz <= 10'd613/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==0/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd2;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==1'd1/*MS*/))  xpc10nz <= 10'd612/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd3]!=0/*MS*/) && !xpc10_stall)  begin 
                               TCCl0_12_V_0 <= 32'd1+TCCl0_12_V_0;
                               TCCl0_12_V_1 <= 32'd4;
                               end 
                              if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==1'd1/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd2;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==2'd2/*MS*/))  xpc10nz <= 10'd611/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==2'd2/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd2;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=2'd3/*MS*/) && 
                      (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd3]!=0/*MS*/))  xpc10nz <= 7'd65/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==0/*MS*/)) 
                       xpc10nz <= 10'd617/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==1'd1/*MS*/)) 
                       xpc10nz <= 10'd616/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==2'd2/*MS*/)) 
                       xpc10nz <= 10'd615/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==2'd3/*MS*/)) 
                       xpc10nz <= 10'd614/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==2'd3/*MS*/))  xpc10nz <= 10'd610/*xpc10nz*/;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==0/*MS*/) && 
                      !xpc10_stall)  TCCl0_12_V_1 <= 32'd3;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==1'd1/*MS*/) && 
                      !xpc10_stall)  TCCl0_12_V_1 <= 32'd3;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==2'd2/*MS*/) && 
                      !xpc10_stall)  TCCl0_12_V_1 <= 32'd3;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd3/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=2'd2/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0
                      [2'd2]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd2]!=0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==2'd3/*MS*/) && 
                      !xpc10_stall)  TCCl0_12_V_1 <= 32'd3;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd2]==2'd3/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd2;
                           end 
                      endcase
              if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==0/*MS*/))  begin if ((xpc10nz==10'd547/*US*/))  xpc10nz <= 10'd548/*xpc10nz*/;
                       end 
                   else if ((xpc10nz==10'd547/*US*/))  xpc10nz <= 7'd65/*xpc10nz*/;
                      
              case (xpc10nz) // synthesis full_case 
                  7'd95/*US*/:  begin 
                      if (!(!TTMT4Main_V_11))  xpc10nz <= 7'd103/*xpc10nz*/;
                           else  xpc10nz <= 7'd96/*xpc10nz*/;
                      if (!(!TTMT4Main_V_11) && !xpc10_stall)  begin 
                               TClo6_9_V_1 <= 32'd0;
                               TTMT4Main_V_13 <= 64'h0;
                               end 
                              if (!TTMT4Main_V_11 && !xpc10_stall)  begin 
                               TTMT4Main_V_13 <= 64'h0;
                               TCl6_SPILL_256 <= -32'd4;
                               end 
                               end 
                      
                  9'd327/*US*/:  begin 
                      if ((A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]==0/*MS*/))  xpc10nz <= 9'd328/*xpc10nz*/;
                           else  xpc10nz <= 9'd323/*xpc10nz*/;
                      if ((A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]==0/*MS*/) && !xpc10_stall)  TCin1_9_V_0 <= TCin1_9_V_6
                          ;

                          if ((A_sA_SINT_CC_SCALbx22_ARB0[A_SINT_CC_SCALbx24_next_victim]!=0/*MS*/) && !xpc10_stall)  begin 
                               TCin1_9_V_2 <= TCin1_9_V_7;
                               TCin1_9_V_0 <= TCin1_9_V_6;
                               end 
                               end 
                      
                  9'd334/*US*/:  begin 
                      if (!(!(32'hffffffff&TCi1_SPILL_256)))  xpc10nz <= 8'd252/*xpc10nz*/;
                           else  xpc10nz <= 8'd251/*xpc10nz*/;
                      if (!(!(32'hffffffff&TCi1_SPILL_256)) && !xpc10_stall)  begin 
                               TTMT4Main_V_7 <= TCi1_SPILL_256;
                               TTMT4Main_V_2 <= 32'd1+TTMT4Main_V_2;
                               end 
                              if (!(32'hffffffff&TCi1_SPILL_256) && !xpc10_stall)  begin 
                               TTMT4Main_V_7 <= TCi1_SPILL_256;
                               TTMT4Main_V_3 <= 32'd1+TTMT4Main_V_3;
                               end 
                               end 
                      
                  9'd338/*US*/:  begin 
                      if ((A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==0/*MS*/))  xpc10nz <= 9'd339/*xpc10nz*/;
                           else  xpc10nz <= 8'd250/*xpc10nz*/;
                      if ((A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]==0/*MS*/) && !xpc10_stall)  TCi1_SPILL_256 <= 32'd0;
                          if ((A_sA_SINT_CC_SCALbx22_ARB0[TCin1_9_V_4]!=0/*MS*/) && !xpc10_stall)  begin 
                               TCi1_SPILL_256 <= 32'd0;
                               TTMT4Main_V_7 <= 32'h0;
                               end 
                               end 
                      
                  10'd534/*US*/:  begin 
                      
                      case (A_sA_SINT_CC_SCALbx20_ARA0[TCCl0_12_V_1]) // synthesis full_case 
                          0/*MS*/:  xpc10nz <= 10'd536/*xpc10nz*/;

                          1'd1/*MS*/:  xpc10nz <= 10'd535/*xpc10nz*/;
                      endcase
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[TCCl0_12_V_1]==1'd1/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd1+TCCl0_12_V_1
                          ;

                          if (((A_sA_SINT_CC_SCALbx20_ARA0[TCCl0_12_V_1]==0/*MS*/)? !xpc10_stall: (A_sA_SINT_CC_SCALbx20_ARA0[TCCl0_12_V_1
                      ]!=1'd1/*MS*/) && !xpc10_stall))  TCCl0_12_V_1 <= 32'd1+TCCl0_12_V_1;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[TCCl0_12_V_1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCCl0_12_V_1]!=0/*MS*/)) 
                       xpc10nz <= 10'd532/*xpc10nz*/;
                           end 
                      
                  10'd547/*US*/:  begin 
                      if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd3]==0/*MS*/) && !xpc10_stall)  TCCl0_12_V_1 <= 32'd4;
                          if ((A_sA_SINT_CC_SCALbx20_ARA0[2'd3]!=0/*MS*/) && !xpc10_stall)  begin 
                               TCCl0_12_V_0 <= 32'd1+TCCl0_12_V_0;
                               TCCl0_12_V_1 <= 32'd4;
                               end 
                               end 
                      endcase
              if ((A_sA_SINT_CC_SCALbx20_ARA0[TCCl0_12_V_1]==0/*MS*/))  begin if ((xpc10nz==10'd537/*US*/))  xpc10nz <= 10'd538/*xpc10nz*/;
                       end 
                   else if ((xpc10nz==10'd537/*US*/))  xpc10nz <= 10'd532/*xpc10nz*/;
                      if (isMODULUS10RRh10vld || isMODULUS10_rdy) 
                  case (xpc10nz) // synthesis full_case 
                      8'd170/*US*/:  xpc10nz <= 8'd236/*xpc10nz*/;

                      8'd235/*US*/:  xpc10nz <= 8'd236/*xpc10nz*/;

                      9'd406/*US*/:  xpc10nz <= 9'd472/*xpc10nz*/;

                      9'd471/*US*/:  xpc10nz <= 9'd472/*xpc10nz*/;
                  endcase
                  if ((TTMT4Main_V_4<15'h_5555)) 
                  case (xpc10nz) // synthesis full_case 
                      7'd86/*US*/:  xpc10nz <= 8'd244/*xpc10nz*/;

                      8'd253/*US*/:  xpc10nz <= 8'd244/*xpc10nz*/;
                  endcase
                   else 
                  case (xpc10nz) // synthesis full_case 
                      7'd86/*US*/:  xpc10nz <= 7'd87/*xpc10nz*/;

                      8'd253/*US*/:  xpc10nz <= 7'd87/*xpc10nz*/;
                  endcase
              if ((TTMT4Main_V_4<15'h_5555) && (xpc10nz==7'd86/*US*/) && !xpc10_stall)  A_SINT_CC_SCALbx28_seed <= 32'h_2aa0_1d31+32'h_7ff8_a3ed
                  *A_SINT_CC_SCALbx28_seed;

                  
              case (xpc10nz) // synthesis full_case 
                  7'd99/*US*/:  begin 
                      if ((TTMT4Main_V_10<15'h_5555))  xpc10nz <= 7'd90/*xpc10nz*/;
                           else  xpc10nz <= 7'd100/*xpc10nz*/;
                      if ((TTMT4Main_V_10<15'h_5555) && !xpc10_stall)  A_SINT_CC_SCALbx28_seed <= 32'h_2aa0_1d31+32'h_7ff8_a3ed*A_SINT_CC_SCALbx28_seed
                          ;

                           end 
                      
                  7'd106/*US*/:  begin 
                      if ((TCha3_10_V_0<0))  xpc10nz <= 8'd171/*xpc10nz*/;
                           else  xpc10nz <= 7'd107/*xpc10nz*/;
                      if ((TCha3_10_V_0<0) && !xpc10_stall)  TCha3_10_V_0 <= (0-TCha3_10_V_0);
                           isMODULUS10RRh10primed <= !xpc10_stall;
                       end 
                      
                  8'd238/*US*/:  begin 
                      if (!TTMT4Main_V_14 && (TTMT4Main_V_12==TTMT4Main_V_13) && !xpc10_stall)  TTMT4Main_V_9 <= 32'd1+TTMT4Main_V_9;
                          if ((!(!TTMT4Main_V_14)? !xpc10_stall: (TTMT4Main_V_12!=TTMT4Main_V_13) && !xpc10_stall))  TTMT4Main_V_8 <= 32'd1
                          +TTMT4Main_V_8;

                          if (!TTMT4Main_V_14 && (TTMT4Main_V_12==TTMT4Main_V_13))  xpc10nz <= 7'd97/*xpc10nz*/;
                          if ((!(!TTMT4Main_V_14)? 1'd1: (TTMT4Main_V_12!=TTMT4Main_V_13)))  xpc10nz <= 7'd98/*xpc10nz*/;
                           end 
                      
                  8'd250/*US*/:  begin 
                      if (!(!TTMT4Main_V_7))  xpc10nz <= 8'd252/*xpc10nz*/;
                           else  xpc10nz <= 8'd251/*xpc10nz*/;
                      if (!TTMT4Main_V_7 && !xpc10_stall)  TTMT4Main_V_3 <= 32'd1+TTMT4Main_V_3;
                          if (!(!TTMT4Main_V_7) && !xpc10_stall)  TTMT4Main_V_2 <= 32'd1+TTMT4Main_V_2;
                           end 
                      endcase
              if ((TTMT4Main_V_4<15'h_5555) && (xpc10nz==8'd253/*US*/) && !xpc10_stall)  A_SINT_CC_SCALbx28_seed <= 32'h_2aa0_1d31+32'h_7ff8_a3ed
                  *A_SINT_CC_SCALbx28_seed;

                  
              case (xpc10nz) // synthesis full_case 
                  7'd100/*US*/:  xpc10nz <= 7'd101/*xpc10nz*/;

                  7'd101/*US*/:  xpc10nz <= 7'd102/*xpc10nz*/;

                  9'd342/*US*/:  begin 
                      if ((TCha6_10_V_0<0))  xpc10nz <= 9'd407/*xpc10nz*/;
                           else  xpc10nz <= 9'd343/*xpc10nz*/;
                      if ((TCha6_10_V_0<0) && !xpc10_stall)  TCha6_10_V_0 <= (0-TCha6_10_V_0);
                           isMODULUS10RRh10primed <= !xpc10_stall;
                       end 
                      
                  10'd532/*US*/:  begin 
                      if ((TCCl0_12_V_1<3'd4))  xpc10nz <= 10'd533/*xpc10nz*/;
                           else  xpc10nz <= 7'd65/*xpc10nz*/;
                      if ((((A_sA_SINT_CC_SCALbx20_ARA0[TCCl0_12_V_1]==2'd3/*MS*/)? 1'd1: (A_sA_SINT_CC_SCALbx20_ARA0[TCCl0_12_V_1]!=
                      0/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCCl0_12_V_1]!=1'd1/*MS*/) && (A_sA_SINT_CC_SCALbx20_ARA0[TCCl0_12_V_1]
                      !=2'd2/*MS*/)) || (A_sA_SINT_CC_SCALbx20_ARA0[TCCl0_12_V_1]==0/*MS*/) || (A_sA_SINT_CC_SCALbx20_ARA0[TCCl0_12_V_1
                      ]==1'd1/*MS*/) || (A_sA_SINT_CC_SCALbx20_ARA0[TCCl0_12_V_1]==2'd2/*MS*/)) && !xpc10_stall && (TCCl0_12_V_1<3'd4
                      ))  TCCl0_12_V_1 <= 32'd1+TCCl0_12_V_1;
                          if ((TCCl0_12_V_1>=3'd4) && !xpc10_stall)  TCCl0_12_V_0 <= 32'd1+TCCl0_12_V_0;
                           end 
                      endcase
              if (isMODULUS10_rdy && isMODULUS10RRh10primed)  begin 
                       isMODULUS10RRh10primed <= 1'd0;
                       isMODULUS10RRh10vld <= 1'd1;
                       isMODULUS10RRh10hold <= isMODULUS10_RR;
                       end 
                      if (SINTCCMAPR12NoCE0ARB0RRh10shot0)  begin 
                       SINTCCMAPR12NoCE0ARB0RRh10hold <= A_SINT_CC_MAPR12NoCE0_ARB0_RDD0;
                       SINTCCMAPR12NoCE0ARB0RRh10hold <= A_SINT_CC_MAPR12NoCE0_ARB0_RDD0;
                       SINTCCMAPR12NoCE0ARB0RRh10hold <= A_SINT_CC_MAPR12NoCE0_ARB0_RDD0;
                       end 
                      if (SINTCCMAPR12NoCE1ARB0RRh10shot0)  begin 
                       SINTCCMAPR12NoCE1ARB0RRh10hold <= A_SINT_CC_MAPR12NoCE1_ARB0_RDD0;
                       SINTCCMAPR12NoCE1ARB0RRh10hold <= A_SINT_CC_MAPR12NoCE1_ARB0_RDD0;
                       SINTCCMAPR12NoCE1ARB0RRh10hold <= A_SINT_CC_MAPR12NoCE1_ARB0_RDD0;
                       end 
                      if (SINTCCMAPR12NoCE2ARB0RRh10shot0)  begin 
                       SINTCCMAPR12NoCE2ARB0RRh10hold <= A_SINT_CC_MAPR12NoCE2_ARB0_RDD0;
                       SINTCCMAPR12NoCE2ARB0RRh10hold <= A_SINT_CC_MAPR12NoCE2_ARB0_RDD0;
                       SINTCCMAPR12NoCE2ARB0RRh10hold <= A_SINT_CC_MAPR12NoCE2_ARB0_RDD0;
                       end 
                      if (SINTCCMAPR12NoCE3ARB0RRh10shot0)  begin 
                       SINTCCMAPR12NoCE3ARB0RRh10hold <= A_SINT_CC_MAPR12NoCE3_ARB0_RDD0;
                       SINTCCMAPR12NoCE3ARB0RRh10hold <= A_SINT_CC_MAPR12NoCE3_ARB0_RDD0;
                       SINTCCMAPR12NoCE3ARB0RRh10hold <= A_SINT_CC_MAPR12NoCE3_ARB0_RDD0;
                       end 
                      if (SINTCCMAPR10NoCE0ARA0RRh10shot0)  begin 
                       SINTCCMAPR10NoCE0ARA0RRh10hold <= A_SINT_CC_MAPR10NoCE0_ARA0_RDD0;
                       SINTCCMAPR10NoCE0ARA0RRh10hold <= A_SINT_CC_MAPR10NoCE0_ARA0_RDD0;
                       SINTCCMAPR10NoCE0ARA0RRh10hold <= A_SINT_CC_MAPR10NoCE0_ARA0_RDD0;
                       end 
                      if (SINTCCMAPR10NoCE1ARA0RRh10shot0)  begin 
                       SINTCCMAPR10NoCE1ARA0RRh10hold <= A_SINT_CC_MAPR10NoCE1_ARA0_RDD0;
                       SINTCCMAPR10NoCE1ARA0RRh10hold <= A_SINT_CC_MAPR10NoCE1_ARA0_RDD0;
                       SINTCCMAPR10NoCE1ARA0RRh10hold <= A_SINT_CC_MAPR10NoCE1_ARA0_RDD0;
                       end 
                      if (SINTCCMAPR10NoCE2ARA0RRh10shot0)  begin 
                       SINTCCMAPR10NoCE2ARA0RRh10hold <= A_SINT_CC_MAPR10NoCE2_ARA0_RDD0;
                       SINTCCMAPR10NoCE2ARA0RRh10hold <= A_SINT_CC_MAPR10NoCE2_ARA0_RDD0;
                       SINTCCMAPR10NoCE2ARA0RRh10hold <= A_SINT_CC_MAPR10NoCE2_ARA0_RDD0;
                       end 
                      if (SINTCCMAPR10NoCE3ARA0RRh10shot0)  begin 
                       SINTCCMAPR10NoCE3ARA0RRh10hold <= A_SINT_CC_MAPR10NoCE3_ARA0_RDD0;
                       SINTCCMAPR10NoCE3ARA0RRh10hold <= A_SINT_CC_MAPR10NoCE3_ARA0_RDD0;
                       SINTCCMAPR10NoCE3ARA0RRh10hold <= A_SINT_CC_MAPR10NoCE3_ARA0_RDD0;
                       end 
                      
              case (xpc10nz) // synthesis full_case 
                  1'd1/*US*/:  xpc10nz <= 2'd2/*US*/;

                  3'd4/*US*/:  xpc10nz <= 3'd5/*xpc10nz*/;

                  3'd5/*US*/:  xpc10nz <= 3'd6/*US*/;

                  3'd7/*US*/:  xpc10nz <= 4'd8/*xpc10nz*/;

                  4'd8/*US*/:  xpc10nz <= 4'd9/*US*/;

                  4'd10/*US*/:  xpc10nz <= 4'd11/*US*/;

                  4'd12/*US*/:  xpc10nz <= 4'd13/*xpc10nz*/;

                  4'd13/*US*/:  xpc10nz <= 4'd14/*US*/;

                  4'd15/*US*/:  xpc10nz <= 5'd16/*xpc10nz*/;

                  5'd16/*US*/:  xpc10nz <= 5'd17/*US*/;

                  5'd19/*US*/:  xpc10nz <= 5'd20/*xpc10nz*/;

                  7'd64/*US*/:  xpc10nz <= 7'd65/*xpc10nz*/;

                  7'd82/*US*/:  xpc10nz <= 7'd83/*xpc10nz*/;

                  7'd83/*US*/:  xpc10nz <= 7'd84/*xpc10nz*/;

                  7'd84/*US*/:  xpc10nz <= 7'd85/*xpc10nz*/;

                  7'd85/*US*/:  xpc10nz <= 7'd86/*xpc10nz*/;

                  7'd87/*US*/:  xpc10nz <= 7'd88/*xpc10nz*/;

                  7'd88/*US*/:  xpc10nz <= 7'd89/*xpc10nz*/;

                  7'd89/*US*/:  xpc10nz <= 7'd90/*xpc10nz*/;

                  7'd90/*US*/:  xpc10nz <= 7'd91/*xpc10nz*/;

                  7'd91/*US*/:  xpc10nz <= 7'd92/*xpc10nz*/;

                  7'd92/*US*/:  xpc10nz <= 7'd93/*xpc10nz*/;

                  7'd93/*US*/:  xpc10nz <= 7'd94/*xpc10nz*/;

                  7'd94/*US*/:  xpc10nz <= 7'd95/*xpc10nz*/;

                  7'd97/*US*/:  xpc10nz <= 7'd98/*xpc10nz*/;

                  7'd98/*US*/:  xpc10nz <= 7'd99/*xpc10nz*/;

                  7'd102/*US*/:  xpc10nz <= 7'd102/*xpc10nz*/;

                  7'd103/*US*/:  xpc10nz <= 7'd104/*xpc10nz*/;

                  7'd104/*US*/:  xpc10nz <= 7'd105/*xpc10nz*/;

                  7'd105/*US*/:  xpc10nz <= 7'd106/*xpc10nz*/;

                  8'd170/*US*/: if ((TCha3_10_V_0>=0) && !xpc10_stall)  TClo6_9_V_1 <= (isMODULUS10RRh10vld? isMODULUS10RRh10hold: isMODULUS10_RR
                      );

                      
                  8'd171/*US*/:  begin 
                       isMODULUS10RRh10primed <= !xpc10_stall;
                       xpc10nz <= 8'd172/*xpc10nz*/;
                       end 
                      
                  8'd240/*US*/:  xpc10nz <= 8'd241/*xpc10nz*/;

                  8'd241/*US*/:  xpc10nz <= 8'd238/*xpc10nz*/;

                  8'd243/*US*/:  begin 
                      if ((TClo6_9_V_0>=3'd4) && (TClo6_9_V_0!=3'd4/*US*/) && !xpc10_stall)  TClo6_9_V_2 <= ((A_sA_SINT_CC_SCALbx22_ARB0
                          [TClo6_9_V_0]==2'd3/*MS*/)? ((xpc10nz==8'd243/*US*/)? A_SINT_CC_MAPR12NoCE3_ARB0_RDD0: SINTCCMAPR12NoCE3ARB0RRh10hold
                          ): ((A_sA_SINT_CC_SCALbx22_ARB0[TClo6_9_V_0]==2'd2/*MS*/)? ((xpc10nz==8'd243/*US*/)? A_SINT_CC_MAPR12NoCE2_ARB0_RDD0
                          : SINTCCMAPR12NoCE2ARB0RRh10hold): ((A_sA_SINT_CC_SCALbx22_ARB0[TClo6_9_V_0]==1'd1/*MS*/)? ((xpc10nz==8'd243
                          /*US*/)? A_SINT_CC_MAPR12NoCE1_ARB0_RDD0: SINTCCMAPR12NoCE1ARB0RRh10hold): ((A_sA_SINT_CC_SCALbx22_ARB0[TClo6_9_V_0
                          ]==0/*MS*/)? ((xpc10nz==8'd243/*US*/)? A_SINT_CC_MAPR12NoCE0_ARB0_RDD0: SINTCCMAPR12NoCE0ARB0RRh10hold): 32'bx
                          ))));

                           xpc10nz <= 8'd239/*xpc10nz*/;
                       end 
                      
                  8'd244/*US*/:  xpc10nz <= 8'd245/*xpc10nz*/;

                  8'd245/*US*/:  xpc10nz <= 8'd246/*xpc10nz*/;

                  8'd246/*US*/:  xpc10nz <= 8'd247/*xpc10nz*/;

                  8'd247/*US*/:  xpc10nz <= 8'd248/*xpc10nz*/;

                  8'd248/*US*/:  xpc10nz <= 8'd249/*xpc10nz*/;

                  8'd251/*US*/:  xpc10nz <= 8'd252/*xpc10nz*/;

                  8'd252/*US*/:  xpc10nz <= 8'd253/*xpc10nz*/;

                  8'd254/*US*/:  xpc10nz <= 8'd255/*xpc10nz*/;

                  8'd255/*US*/:  xpc10nz <= 9'd256/*xpc10nz*/;

                  9'd257/*US*/:  xpc10nz <= 9'd258/*xpc10nz*/;

                  9'd258/*US*/:  xpc10nz <= 9'd259/*xpc10nz*/;

                  9'd284/*US*/:  xpc10nz <= 9'd285/*xpc10nz*/;

                  9'd286/*US*/:  xpc10nz <= 9'd287/*xpc10nz*/;

                  9'd288/*US*/:  xpc10nz <= 9'd289/*xpc10nz*/;

                  9'd318/*US*/:  xpc10nz <= 9'd319/*xpc10nz*/;

                  9'd319/*US*/:  xpc10nz <= 9'd320/*xpc10nz*/;

                  9'd320/*US*/:  xpc10nz <= 9'd321/*xpc10nz*/;

                  9'd321/*US*/:  xpc10nz <= 9'd322/*xpc10nz*/;

                  9'd322/*US*/:  xpc10nz <= 9'd259/*xpc10nz*/;

                  9'd323/*US*/:  xpc10nz <= 9'd320/*xpc10nz*/;

                  9'd329/*US*/:  xpc10nz <= 9'd323/*xpc10nz*/;

                  9'd340/*US*/:  xpc10nz <= 8'd250/*xpc10nz*/;

                  9'd341/*US*/:  xpc10nz <= 9'd342/*xpc10nz*/;

                  9'd406/*US*/: if ((TCha6_10_V_0>=0) && !xpc10_stall)  TCin1_9_V_5 <= (isMODULUS10RRh10vld? isMODULUS10RRh10hold: isMODULUS10_RR
                      );

                      
                  9'd407/*US*/:  begin 
                       isMODULUS10RRh10primed <= !xpc10_stall;
                       xpc10nz <= 9'd408/*xpc10nz*/;
                       end 
                      
                  9'd502/*US*/:  xpc10nz <= 9'd284/*xpc10nz*/;

                  10'd539/*US*/:  xpc10nz <= 10'd532/*xpc10nz*/;

                  10'd549/*US*/:  xpc10nz <= 7'd65/*xpc10nz*/;
              endcase
              if (Z64USCCSCALbx26ARA0RRh10shot0)  Z64USCCSCALbx26ARA0RRh10hold <= A_64_US_CC_SCALbx26_ARA0_RDD0;
                  if (!xpc10_stall && xpc10_clear)  isMODULUS10RRh10vld <= 1'd0;
                   SINTCCMAPR10NoCE0ARA0RRh10shot0 <= ((xpc10nz==9'd472/*US*/) || (xpc10nz==8'd236/*US*/) || (xpc10nz==9'd285/*US*/)) && 
              !xpc10_stall;

               SINTCCMAPR10NoCE1ARA0RRh10shot0 <= ((xpc10nz==9'd472/*US*/) || (xpc10nz==8'd236/*US*/) || (xpc10nz==9'd285/*US*/)) && 
              !xpc10_stall;

               SINTCCMAPR10NoCE2ARA0RRh10shot0 <= ((xpc10nz==9'd472/*US*/) || (xpc10nz==8'd236/*US*/) || (xpc10nz==9'd285/*US*/)) && 
              !xpc10_stall;

               SINTCCMAPR10NoCE3ARA0RRh10shot0 <= ((xpc10nz==9'd472/*US*/) || (xpc10nz==8'd236/*US*/) || (xpc10nz==9'd285/*US*/)) && 
              !xpc10_stall;

               SINTCCMAPR12NoCE0ARB0RRh10shot0 <= (((TClo6_9_V_0>=3'd4) && (xpc10nz==8'd242/*US*/) || (xpc10nz==8'd236/*US*/) && (TTMT4Main_V_11
              ==((A_sA_SINT_CC_SCALbx20_ARA0[TClo6_9_V_0]==2'd3/*MS*/)? ((xpc10nz==8'd237/*US*/)? A_SINT_CC_MAPR10NoCE3_ARA0_RDD0: SINTCCMAPR10NoCE3ARA0RRh10hold
              ): ((A_sA_SINT_CC_SCALbx20_ARA0[TClo6_9_V_0]==2'd2/*MS*/)? ((xpc10nz==8'd237/*US*/)? A_SINT_CC_MAPR10NoCE2_ARA0_RDD0: SINTCCMAPR10NoCE2ARA0RRh10hold
              ): ((A_sA_SINT_CC_SCALbx20_ARA0[TClo6_9_V_0]==1'd1/*MS*/)? ((xpc10nz==8'd237/*US*/)? A_SINT_CC_MAPR10NoCE1_ARA0_RDD0: SINTCCMAPR10NoCE1ARA0RRh10hold
              ): ((A_sA_SINT_CC_SCALbx20_ARA0[TClo6_9_V_0]==0/*MS*/)? ((xpc10nz==8'd237/*US*/)? A_SINT_CC_MAPR10NoCE0_ARA0_RDD0: SINTCCMAPR10NoCE0ARA0RRh10hold
              ): 1'bx)))))) && (TClo6_9_V_0!=3'd4/*US*/) || (xpc10nz==9'd287/*US*/)) && !xpc10_stall;

               SINTCCMAPR12NoCE1ARB0RRh10shot0 <= (((TClo6_9_V_0>=3'd4) && (xpc10nz==8'd242/*US*/) || (xpc10nz==8'd236/*US*/) && (TTMT4Main_V_11
              ==((A_sA_SINT_CC_SCALbx20_ARA0[TClo6_9_V_0]==2'd3/*MS*/)? ((xpc10nz==8'd237/*US*/)? A_SINT_CC_MAPR10NoCE3_ARA0_RDD0: SINTCCMAPR10NoCE3ARA0RRh10hold
              ): ((A_sA_SINT_CC_SCALbx20_ARA0[TClo6_9_V_0]==2'd2/*MS*/)? ((xpc10nz==8'd237/*US*/)? A_SINT_CC_MAPR10NoCE2_ARA0_RDD0: SINTCCMAPR10NoCE2ARA0RRh10hold
              ): ((A_sA_SINT_CC_SCALbx20_ARA0[TClo6_9_V_0]==1'd1/*MS*/)? ((xpc10nz==8'd237/*US*/)? A_SINT_CC_MAPR10NoCE1_ARA0_RDD0: SINTCCMAPR10NoCE1ARA0RRh10hold
              ): ((A_sA_SINT_CC_SCALbx20_ARA0[TClo6_9_V_0]==0/*MS*/)? ((xpc10nz==8'd237/*US*/)? A_SINT_CC_MAPR10NoCE0_ARA0_RDD0: SINTCCMAPR10NoCE0ARA0RRh10hold
              ): 1'bx)))))) && (TClo6_9_V_0!=3'd4/*US*/) || (xpc10nz==9'd287/*US*/)) && !xpc10_stall;

               SINTCCMAPR12NoCE2ARB0RRh10shot0 <= (((TClo6_9_V_0>=3'd4) && (xpc10nz==8'd242/*US*/) || (xpc10nz==8'd236/*US*/) && (TTMT4Main_V_11
              ==((A_sA_SINT_CC_SCALbx20_ARA0[TClo6_9_V_0]==2'd3/*MS*/)? ((xpc10nz==8'd237/*US*/)? A_SINT_CC_MAPR10NoCE3_ARA0_RDD0: SINTCCMAPR10NoCE3ARA0RRh10hold
              ): ((A_sA_SINT_CC_SCALbx20_ARA0[TClo6_9_V_0]==2'd2/*MS*/)? ((xpc10nz==8'd237/*US*/)? A_SINT_CC_MAPR10NoCE2_ARA0_RDD0: SINTCCMAPR10NoCE2ARA0RRh10hold
              ): ((A_sA_SINT_CC_SCALbx20_ARA0[TClo6_9_V_0]==1'd1/*MS*/)? ((xpc10nz==8'd237/*US*/)? A_SINT_CC_MAPR10NoCE1_ARA0_RDD0: SINTCCMAPR10NoCE1ARA0RRh10hold
              ): ((A_sA_SINT_CC_SCALbx20_ARA0[TClo6_9_V_0]==0/*MS*/)? ((xpc10nz==8'd237/*US*/)? A_SINT_CC_MAPR10NoCE0_ARA0_RDD0: SINTCCMAPR10NoCE0ARA0RRh10hold
              ): 1'bx)))))) && (TClo6_9_V_0!=3'd4/*US*/) || (xpc10nz==9'd287/*US*/)) && !xpc10_stall;

               SINTCCMAPR12NoCE3ARB0RRh10shot0 <= (((TClo6_9_V_0>=3'd4) && (xpc10nz==8'd242/*US*/) || (xpc10nz==8'd236/*US*/) && (TTMT4Main_V_11
              ==((A_sA_SINT_CC_SCALbx20_ARA0[TClo6_9_V_0]==2'd3/*MS*/)? ((xpc10nz==8'd237/*US*/)? A_SINT_CC_MAPR10NoCE3_ARA0_RDD0: SINTCCMAPR10NoCE3ARA0RRh10hold
              ): ((A_sA_SINT_CC_SCALbx20_ARA0[TClo6_9_V_0]==2'd2/*MS*/)? ((xpc10nz==8'd237/*US*/)? A_SINT_CC_MAPR10NoCE2_ARA0_RDD0: SINTCCMAPR10NoCE2ARA0RRh10hold
              ): ((A_sA_SINT_CC_SCALbx20_ARA0[TClo6_9_V_0]==1'd1/*MS*/)? ((xpc10nz==8'd237/*US*/)? A_SINT_CC_MAPR10NoCE1_ARA0_RDD0: SINTCCMAPR10NoCE1ARA0RRh10hold
              ): ((A_sA_SINT_CC_SCALbx20_ARA0[TClo6_9_V_0]==0/*MS*/)? ((xpc10nz==8'd237/*US*/)? A_SINT_CC_MAPR10NoCE0_ARA0_RDD0: SINTCCMAPR10NoCE0ARA0RRh10hold
              ): 1'bx)))))) && (TClo6_9_V_0!=3'd4/*US*/) || (xpc10nz==9'd287/*US*/)) && !xpc10_stall;

               Z64USCCSCALbx26ARA0RRh10shot0 <= (xpc10nz==8'd239/*US*/) && !xpc10_stall;
               xpc10_trk64 <= ((7'd64/*MS*/==-11'd609+xpc10nz) || (7'd64/*MS*/==-11'd599+xpc10nz) || (7'd64/*MS*/==-11'd588+xpc10nz) || 
              (7'd64/*MS*/==-11'd576+xpc10nz) || (7'd64/*MS*/==-11'd571+xpc10nz) || (7'd64/*MS*/==-11'd565+xpc10nz) || (7'd64/*MS*/==
              -11'd558+xpc10nz) || (7'd64/*MS*/==-11'd550+xpc10nz) || (7'd64/*MS*/==-11'd549+xpc10nz) || (7'd64/*MS*/==-11'd547+xpc10nz
              ) || (7'd64/*MS*/==-11'd544+xpc10nz) || (7'd64/*MS*/==-11'd540+xpc10nz) || (7'd64/*MS*/==-11'd539+xpc10nz) || (7'd64/*MS*/==
              -11'd537+xpc10nz) || (7'd64/*MS*/==-11'd534+xpc10nz) || (7'd64/*MS*/==-11'd532+xpc10nz) || (7'd64/*MS*/==-11'd528+xpc10nz
              ) || (7'd64/*MS*/==-10'd503+xpc10nz) || (7'd64/*MS*/==-10'd502+xpc10nz) || (7'd64/*MS*/==-10'd472+xpc10nz) || (7'd64/*MS*/==
              -10'd407+xpc10nz) || (7'd64/*MS*/==-10'd342+xpc10nz) || (7'd64/*MS*/==-10'd341+xpc10nz) || (7'd64/*MS*/==-10'd340+xpc10nz
              ) || (7'd64/*MS*/==-10'd338+xpc10nz) || (7'd64/*MS*/==-10'd335+xpc10nz) || (7'd64/*MS*/==-10'd334+xpc10nz) || (7'd64/*MS*/==
              -10'd330+xpc10nz) || (7'd64/*MS*/==-10'd329+xpc10nz) || (7'd64/*MS*/==-10'd327+xpc10nz) || (7'd64/*MS*/==-10'd324+xpc10nz
              ) || (7'd64/*MS*/==-10'd323+xpc10nz) || (7'd64/*MS*/==-10'd322+xpc10nz) || (7'd64/*MS*/==-10'd321+xpc10nz) || (7'd64/*MS*/==
              -10'd320+xpc10nz) || (7'd64/*MS*/==-10'd319+xpc10nz) || (7'd64/*MS*/==-10'd318+xpc10nz) || (7'd64/*MS*/==-10'd314+xpc10nz
              ) || (7'd64/*MS*/==-10'd289+xpc10nz) || (7'd64/*MS*/==-10'd287+xpc10nz) || (7'd64/*MS*/==-10'd285+xpc10nz) || (7'd64/*MS*/==
              -10'd284+xpc10nz) || (7'd64/*MS*/==-10'd259+xpc10nz) || (7'd64/*MS*/==-10'd258+xpc10nz) || (7'd64/*MS*/==-10'd257+xpc10nz
              ) || (7'd64/*MS*/==-9'd255+xpc10nz) || (7'd64/*MS*/==-9'd254+xpc10nz) || (7'd64/*MS*/==-9'd253+xpc10nz) || (7'd64/*MS*/==
              -9'd252+xpc10nz) || (7'd64/*MS*/==-9'd251+xpc10nz) || (7'd64/*MS*/==-9'd250+xpc10nz) || (7'd64/*MS*/==-9'd249+xpc10nz) || 
              (7'd64/*MS*/==-9'd248+xpc10nz) || (7'd64/*MS*/==-9'd247+xpc10nz) || (7'd64/*MS*/==-9'd246+xpc10nz) || (7'd64/*MS*/==-9'd245
              +xpc10nz) || (7'd64/*MS*/==-9'd244+xpc10nz) || (7'd64/*MS*/==-9'd242+xpc10nz) || (7'd64/*MS*/==-9'd241+xpc10nz) || (7'd64
              /*MS*/==-9'd239+xpc10nz) || (7'd64/*MS*/==-9'd238+xpc10nz) || (7'd64/*MS*/==-9'd236+xpc10nz) || (7'd64/*MS*/==-9'd171+xpc10nz
              ) || (7'd64/*MS*/==-8'd106+xpc10nz) || (7'd64/*MS*/==-8'd105+xpc10nz) || (7'd64/*MS*/==-8'd104+xpc10nz) || (7'd64/*MS*/==
              -8'd103+xpc10nz) || (7'd64/*MS*/==-8'd102+xpc10nz) || (7'd64/*MS*/==-8'd101+xpc10nz) || (7'd64/*MS*/==-8'd100+xpc10nz) || 
              (7'd64/*MS*/==-8'd99+xpc10nz) || (7'd64/*MS*/==-8'd98+xpc10nz) || (7'd64/*MS*/==-8'd97+xpc10nz) || (7'd64/*MS*/==-8'd96
              +xpc10nz) || (7'd64/*MS*/==-8'd95+xpc10nz) || (7'd64/*MS*/==-8'd94+xpc10nz) || (7'd64/*MS*/==-8'd93+xpc10nz) || (7'd64/*MS*/==
              -8'd92+xpc10nz) || (7'd64/*MS*/==-8'd91+xpc10nz) || (7'd64/*MS*/==-8'd90+xpc10nz) || (7'd64/*MS*/==-8'd89+xpc10nz) || (7'd64
              /*MS*/==-8'd88+xpc10nz) || (7'd64/*MS*/==-8'd87+xpc10nz) || (7'd64/*MS*/==-8'd86+xpc10nz) || (7'd64/*MS*/==-8'd85+xpc10nz
              ) || (7'd64/*MS*/==-8'd84+xpc10nz) || (7'd64/*MS*/==-8'd83+xpc10nz) || (7'd64/*MS*/==-8'd82+xpc10nz) || (7'd64/*MS*/==-8'd65
              +xpc10nz) || (7'd64/*MS*/==-8'd64+xpc10nz) || (7'd64/*MS*/==-7'd59+xpc10nz) || (7'd64/*MS*/==-7'd50+xpc10nz) || (7'd64/*MS*/==
              -7'd37+xpc10nz) || (7'd64/*MS*/==-6'd20+xpc10nz) || (7'd64/*MS*/==-6'd19+xpc10nz) || (7'd64/*MS*/==-6'd18+xpc10nz) || (7'd64
              /*MS*/==-6'd17+xpc10nz) || (7'd64/*MS*/==-6'd16+xpc10nz) || (7'd64/*MS*/==-5'd15+xpc10nz) || (7'd64/*MS*/==-5'd14+xpc10nz
              ) || (7'd64/*MS*/==-5'd13+xpc10nz) || (7'd64/*MS*/==-5'd12+xpc10nz) || (7'd64/*MS*/==-5'd11+xpc10nz) || (7'd64/*MS*/==-5'd10
              +xpc10nz) || (7'd64/*MS*/==-5'd9+xpc10nz) || (7'd64/*MS*/==-5'd8+xpc10nz) || (7'd64/*MS*/==-4'd7+xpc10nz) || (7'd64/*MS*/==
              -4'd6+xpc10nz) || (7'd64/*MS*/==-4'd5+xpc10nz) || (7'd64/*MS*/==-4'd4+xpc10nz) || (7'd64/*MS*/==-3'd3+xpc10nz) || (7'd64
              /*MS*/==-3'd2+xpc10nz) || (7'd64/*MS*/==-2'd1+xpc10nz) || (xpc10nz==7'd64/*US*/)) && !xpc10_clear && !xpc10_stall;

               xpc10_trk63 <= ((6'd63/*MS*/==-11'd609+xpc10nz) || (6'd63/*MS*/==-11'd599+xpc10nz) || (6'd63/*MS*/==-11'd588+xpc10nz) || 
              (6'd63/*MS*/==-11'd576+xpc10nz) || (6'd63/*MS*/==-11'd571+xpc10nz) || (6'd63/*MS*/==-11'd565+xpc10nz) || (6'd63/*MS*/==
              -11'd558+xpc10nz) || (6'd63/*MS*/==-11'd550+xpc10nz) || (6'd63/*MS*/==-11'd549+xpc10nz) || (6'd63/*MS*/==-11'd547+xpc10nz
              ) || (6'd63/*MS*/==-11'd544+xpc10nz) || (6'd63/*MS*/==-11'd540+xpc10nz) || (6'd63/*MS*/==-11'd539+xpc10nz) || (6'd63/*MS*/==
              -11'd537+xpc10nz) || (6'd63/*MS*/==-11'd534+xpc10nz) || (6'd63/*MS*/==-11'd532+xpc10nz) || (6'd63/*MS*/==-11'd528+xpc10nz
              ) || (6'd63/*MS*/==-10'd503+xpc10nz) || (6'd63/*MS*/==-10'd502+xpc10nz) || (6'd63/*MS*/==-10'd472+xpc10nz) || (6'd63/*MS*/==
              -10'd407+xpc10nz) || (6'd63/*MS*/==-10'd342+xpc10nz) || (6'd63/*MS*/==-10'd341+xpc10nz) || (6'd63/*MS*/==-10'd340+xpc10nz
              ) || (6'd63/*MS*/==-10'd338+xpc10nz) || (6'd63/*MS*/==-10'd335+xpc10nz) || (6'd63/*MS*/==-10'd334+xpc10nz) || (6'd63/*MS*/==
              -10'd330+xpc10nz) || (6'd63/*MS*/==-10'd329+xpc10nz) || (6'd63/*MS*/==-10'd327+xpc10nz) || (6'd63/*MS*/==-10'd324+xpc10nz
              ) || (6'd63/*MS*/==-10'd323+xpc10nz) || (6'd63/*MS*/==-10'd322+xpc10nz) || (6'd63/*MS*/==-10'd321+xpc10nz) || (6'd63/*MS*/==
              -10'd320+xpc10nz) || (6'd63/*MS*/==-10'd319+xpc10nz) || (6'd63/*MS*/==-10'd318+xpc10nz) || (6'd63/*MS*/==-10'd314+xpc10nz
              ) || (6'd63/*MS*/==-10'd289+xpc10nz) || (6'd63/*MS*/==-10'd287+xpc10nz) || (6'd63/*MS*/==-10'd285+xpc10nz) || (6'd63/*MS*/==
              -10'd284+xpc10nz) || (6'd63/*MS*/==-10'd259+xpc10nz) || (6'd63/*MS*/==-10'd258+xpc10nz) || (6'd63/*MS*/==-10'd257+xpc10nz
              ) || (6'd63/*MS*/==-9'd255+xpc10nz) || (6'd63/*MS*/==-9'd254+xpc10nz) || (6'd63/*MS*/==-9'd253+xpc10nz) || (6'd63/*MS*/==
              -9'd252+xpc10nz) || (6'd63/*MS*/==-9'd251+xpc10nz) || (6'd63/*MS*/==-9'd250+xpc10nz) || (6'd63/*MS*/==-9'd249+xpc10nz) || 
              (6'd63/*MS*/==-9'd248+xpc10nz) || (6'd63/*MS*/==-9'd247+xpc10nz) || (6'd63/*MS*/==-9'd246+xpc10nz) || (6'd63/*MS*/==-9'd245
              +xpc10nz) || (6'd63/*MS*/==-9'd244+xpc10nz) || (6'd63/*MS*/==-9'd242+xpc10nz) || (6'd63/*MS*/==-9'd241+xpc10nz) || (6'd63
              /*MS*/==-9'd239+xpc10nz) || (6'd63/*MS*/==-9'd238+xpc10nz) || (6'd63/*MS*/==-9'd236+xpc10nz) || (6'd63/*MS*/==-9'd171+xpc10nz
              ) || (6'd63/*MS*/==-8'd106+xpc10nz) || (6'd63/*MS*/==-8'd105+xpc10nz) || (6'd63/*MS*/==-8'd104+xpc10nz) || (6'd63/*MS*/==
              -8'd103+xpc10nz) || (6'd63/*MS*/==-8'd102+xpc10nz) || (6'd63/*MS*/==-8'd101+xpc10nz) || (6'd63/*MS*/==-8'd100+xpc10nz) || 
              (6'd63/*MS*/==-8'd99+xpc10nz) || (6'd63/*MS*/==-8'd98+xpc10nz) || (6'd63/*MS*/==-8'd97+xpc10nz) || (6'd63/*MS*/==-8'd96
              +xpc10nz) || (6'd63/*MS*/==-8'd95+xpc10nz) || (6'd63/*MS*/==-8'd94+xpc10nz) || (6'd63/*MS*/==-8'd93+xpc10nz) || (6'd63/*MS*/==
              -8'd92+xpc10nz) || (6'd63/*MS*/==-8'd91+xpc10nz) || (6'd63/*MS*/==-8'd90+xpc10nz) || (6'd63/*MS*/==-8'd89+xpc10nz) || (6'd63
              /*MS*/==-8'd88+xpc10nz) || (6'd63/*MS*/==-8'd87+xpc10nz) || (6'd63/*MS*/==-8'd86+xpc10nz) || (6'd63/*MS*/==-8'd85+xpc10nz
              ) || (6'd63/*MS*/==-8'd84+xpc10nz) || (6'd63/*MS*/==-8'd83+xpc10nz) || (6'd63/*MS*/==-8'd82+xpc10nz) || (6'd63/*MS*/==-8'd65
              +xpc10nz) || (6'd63/*MS*/==-8'd64+xpc10nz) || (6'd63/*MS*/==-7'd59+xpc10nz) || (6'd63/*MS*/==-7'd50+xpc10nz) || (6'd63/*MS*/==
              -7'd37+xpc10nz) || (6'd63/*MS*/==-6'd20+xpc10nz) || (6'd63/*MS*/==-6'd19+xpc10nz) || (6'd63/*MS*/==-6'd18+xpc10nz) || (6'd63
              /*MS*/==-6'd17+xpc10nz) || (6'd63/*MS*/==-6'd16+xpc10nz) || (6'd63/*MS*/==-5'd15+xpc10nz) || (6'd63/*MS*/==-5'd14+xpc10nz
              ) || (6'd63/*MS*/==-5'd13+xpc10nz) || (6'd63/*MS*/==-5'd12+xpc10nz) || (6'd63/*MS*/==-5'd11+xpc10nz) || (6'd63/*MS*/==-5'd10
              +xpc10nz) || (6'd63/*MS*/==-5'd9+xpc10nz) || (6'd63/*MS*/==-5'd8+xpc10nz) || (6'd63/*MS*/==-4'd7+xpc10nz) || (6'd63/*MS*/==
              -4'd6+xpc10nz) || (6'd63/*MS*/==-4'd5+xpc10nz) || (6'd63/*MS*/==-4'd4+xpc10nz) || (6'd63/*MS*/==-3'd3+xpc10nz) || (6'd63
              /*MS*/==-3'd2+xpc10nz) || (6'd63/*MS*/==-2'd1+xpc10nz) || (xpc10nz==6'd63/*US*/)) && !xpc10_clear && !xpc10_stall;

               xpc10_trk62 <= ((6'd62/*MS*/==-11'd609+xpc10nz) || (6'd62/*MS*/==-11'd599+xpc10nz) || (6'd62/*MS*/==-11'd588+xpc10nz) || 
              (6'd62/*MS*/==-11'd576+xpc10nz) || (6'd62/*MS*/==-11'd571+xpc10nz) || (6'd62/*MS*/==-11'd565+xpc10nz) || (6'd62/*MS*/==
              -11'd558+xpc10nz) || (6'd62/*MS*/==-11'd550+xpc10nz) || (6'd62/*MS*/==-11'd549+xpc10nz) || (6'd62/*MS*/==-11'd547+xpc10nz
              ) || (6'd62/*MS*/==-11'd544+xpc10nz) || (6'd62/*MS*/==-11'd540+xpc10nz) || (6'd62/*MS*/==-11'd539+xpc10nz) || (6'd62/*MS*/==
              -11'd537+xpc10nz) || (6'd62/*MS*/==-11'd534+xpc10nz) || (6'd62/*MS*/==-11'd532+xpc10nz) || (6'd62/*MS*/==-11'd528+xpc10nz
              ) || (6'd62/*MS*/==-10'd503+xpc10nz) || (6'd62/*MS*/==-10'd502+xpc10nz) || (6'd62/*MS*/==-10'd472+xpc10nz) || (6'd62/*MS*/==
              -10'd407+xpc10nz) || (6'd62/*MS*/==-10'd342+xpc10nz) || (6'd62/*MS*/==-10'd341+xpc10nz) || (6'd62/*MS*/==-10'd340+xpc10nz
              ) || (6'd62/*MS*/==-10'd338+xpc10nz) || (6'd62/*MS*/==-10'd335+xpc10nz) || (6'd62/*MS*/==-10'd334+xpc10nz) || (6'd62/*MS*/==
              -10'd330+xpc10nz) || (6'd62/*MS*/==-10'd329+xpc10nz) || (6'd62/*MS*/==-10'd327+xpc10nz) || (6'd62/*MS*/==-10'd324+xpc10nz
              ) || (6'd62/*MS*/==-10'd323+xpc10nz) || (6'd62/*MS*/==-10'd322+xpc10nz) || (6'd62/*MS*/==-10'd321+xpc10nz) || (6'd62/*MS*/==
              -10'd320+xpc10nz) || (6'd62/*MS*/==-10'd319+xpc10nz) || (6'd62/*MS*/==-10'd318+xpc10nz) || (6'd62/*MS*/==-10'd314+xpc10nz
              ) || (6'd62/*MS*/==-10'd289+xpc10nz) || (6'd62/*MS*/==-10'd287+xpc10nz) || (6'd62/*MS*/==-10'd285+xpc10nz) || (6'd62/*MS*/==
              -10'd284+xpc10nz) || (6'd62/*MS*/==-10'd259+xpc10nz) || (6'd62/*MS*/==-10'd258+xpc10nz) || (6'd62/*MS*/==-10'd257+xpc10nz
              ) || (6'd62/*MS*/==-9'd255+xpc10nz) || (6'd62/*MS*/==-9'd254+xpc10nz) || (6'd62/*MS*/==-9'd253+xpc10nz) || (6'd62/*MS*/==
              -9'd252+xpc10nz) || (6'd62/*MS*/==-9'd251+xpc10nz) || (6'd62/*MS*/==-9'd250+xpc10nz) || (6'd62/*MS*/==-9'd249+xpc10nz) || 
              (6'd62/*MS*/==-9'd248+xpc10nz) || (6'd62/*MS*/==-9'd247+xpc10nz) || (6'd62/*MS*/==-9'd246+xpc10nz) || (6'd62/*MS*/==-9'd245
              +xpc10nz) || (6'd62/*MS*/==-9'd244+xpc10nz) || (6'd62/*MS*/==-9'd242+xpc10nz) || (6'd62/*MS*/==-9'd241+xpc10nz) || (6'd62
              /*MS*/==-9'd239+xpc10nz) || (6'd62/*MS*/==-9'd238+xpc10nz) || (6'd62/*MS*/==-9'd236+xpc10nz) || (6'd62/*MS*/==-9'd171+xpc10nz
              ) || (6'd62/*MS*/==-8'd106+xpc10nz) || (6'd62/*MS*/==-8'd105+xpc10nz) || (6'd62/*MS*/==-8'd104+xpc10nz) || (6'd62/*MS*/==
              -8'd103+xpc10nz) || (6'd62/*MS*/==-8'd102+xpc10nz) || (6'd62/*MS*/==-8'd101+xpc10nz) || (6'd62/*MS*/==-8'd100+xpc10nz) || 
              (6'd62/*MS*/==-8'd99+xpc10nz) || (6'd62/*MS*/==-8'd98+xpc10nz) || (6'd62/*MS*/==-8'd97+xpc10nz) || (6'd62/*MS*/==-8'd96
              +xpc10nz) || (6'd62/*MS*/==-8'd95+xpc10nz) || (6'd62/*MS*/==-8'd94+xpc10nz) || (6'd62/*MS*/==-8'd93+xpc10nz) || (6'd62/*MS*/==
              -8'd92+xpc10nz) || (6'd62/*MS*/==-8'd91+xpc10nz) || (6'd62/*MS*/==-8'd90+xpc10nz) || (6'd62/*MS*/==-8'd89+xpc10nz) || (6'd62
              /*MS*/==-8'd88+xpc10nz) || (6'd62/*MS*/==-8'd87+xpc10nz) || (6'd62/*MS*/==-8'd86+xpc10nz) || (6'd62/*MS*/==-8'd85+xpc10nz
              ) || (6'd62/*MS*/==-8'd84+xpc10nz) || (6'd62/*MS*/==-8'd83+xpc10nz) || (6'd62/*MS*/==-8'd82+xpc10nz) || (6'd62/*MS*/==-8'd65
              +xpc10nz) || (6'd62/*MS*/==-8'd64+xpc10nz) || (6'd62/*MS*/==-7'd59+xpc10nz) || (6'd62/*MS*/==-7'd50+xpc10nz) || (6'd62/*MS*/==
              -7'd37+xpc10nz) || (6'd62/*MS*/==-6'd20+xpc10nz) || (6'd62/*MS*/==-6'd19+xpc10nz) || (6'd62/*MS*/==-6'd18+xpc10nz) || (6'd62
              /*MS*/==-6'd17+xpc10nz) || (6'd62/*MS*/==-6'd16+xpc10nz) || (6'd62/*MS*/==-5'd15+xpc10nz) || (6'd62/*MS*/==-5'd14+xpc10nz
              ) || (6'd62/*MS*/==-5'd13+xpc10nz) || (6'd62/*MS*/==-5'd12+xpc10nz) || (6'd62/*MS*/==-5'd11+xpc10nz) || (6'd62/*MS*/==-5'd10
              +xpc10nz) || (6'd62/*MS*/==-5'd9+xpc10nz) || (6'd62/*MS*/==-5'd8+xpc10nz) || (6'd62/*MS*/==-4'd7+xpc10nz) || (6'd62/*MS*/==
              -4'd6+xpc10nz) || (6'd62/*MS*/==-4'd5+xpc10nz) || (6'd62/*MS*/==-4'd4+xpc10nz) || (6'd62/*MS*/==-3'd3+xpc10nz) || (6'd62
              /*MS*/==-3'd2+xpc10nz) || (6'd62/*MS*/==-2'd1+xpc10nz) || (xpc10nz==6'd62/*US*/)) && !xpc10_clear && !xpc10_stall;

               xpc10_trk61 <= ((6'd61/*MS*/==-11'd609+xpc10nz) || (6'd61/*MS*/==-11'd599+xpc10nz) || (6'd61/*MS*/==-11'd588+xpc10nz) || 
              (6'd61/*MS*/==-11'd576+xpc10nz) || (6'd61/*MS*/==-11'd571+xpc10nz) || (6'd61/*MS*/==-11'd565+xpc10nz) || (6'd61/*MS*/==
              -11'd558+xpc10nz) || (6'd61/*MS*/==-11'd550+xpc10nz) || (6'd61/*MS*/==-11'd549+xpc10nz) || (6'd61/*MS*/==-11'd547+xpc10nz
              ) || (6'd61/*MS*/==-11'd544+xpc10nz) || (6'd61/*MS*/==-11'd540+xpc10nz) || (6'd61/*MS*/==-11'd539+xpc10nz) || (6'd61/*MS*/==
              -11'd537+xpc10nz) || (6'd61/*MS*/==-11'd534+xpc10nz) || (6'd61/*MS*/==-11'd532+xpc10nz) || (6'd61/*MS*/==-11'd528+xpc10nz
              ) || (6'd61/*MS*/==-10'd503+xpc10nz) || (6'd61/*MS*/==-10'd502+xpc10nz) || (6'd61/*MS*/==-10'd472+xpc10nz) || (6'd61/*MS*/==
              -10'd407+xpc10nz) || (6'd61/*MS*/==-10'd342+xpc10nz) || (6'd61/*MS*/==-10'd341+xpc10nz) || (6'd61/*MS*/==-10'd340+xpc10nz
              ) || (6'd61/*MS*/==-10'd338+xpc10nz) || (6'd61/*MS*/==-10'd335+xpc10nz) || (6'd61/*MS*/==-10'd334+xpc10nz) || (6'd61/*MS*/==
              -10'd330+xpc10nz) || (6'd61/*MS*/==-10'd329+xpc10nz) || (6'd61/*MS*/==-10'd327+xpc10nz) || (6'd61/*MS*/==-10'd324+xpc10nz
              ) || (6'd61/*MS*/==-10'd323+xpc10nz) || (6'd61/*MS*/==-10'd322+xpc10nz) || (6'd61/*MS*/==-10'd321+xpc10nz) || (6'd61/*MS*/==
              -10'd320+xpc10nz) || (6'd61/*MS*/==-10'd319+xpc10nz) || (6'd61/*MS*/==-10'd318+xpc10nz) || (6'd61/*MS*/==-10'd314+xpc10nz
              ) || (6'd61/*MS*/==-10'd289+xpc10nz) || (6'd61/*MS*/==-10'd287+xpc10nz) || (6'd61/*MS*/==-10'd285+xpc10nz) || (6'd61/*MS*/==
              -10'd284+xpc10nz) || (6'd61/*MS*/==-10'd259+xpc10nz) || (6'd61/*MS*/==-10'd258+xpc10nz) || (6'd61/*MS*/==-10'd257+xpc10nz
              ) || (6'd61/*MS*/==-9'd255+xpc10nz) || (6'd61/*MS*/==-9'd254+xpc10nz) || (6'd61/*MS*/==-9'd253+xpc10nz) || (6'd61/*MS*/==
              -9'd252+xpc10nz) || (6'd61/*MS*/==-9'd251+xpc10nz) || (6'd61/*MS*/==-9'd250+xpc10nz) || (6'd61/*MS*/==-9'd249+xpc10nz) || 
              (6'd61/*MS*/==-9'd248+xpc10nz) || (6'd61/*MS*/==-9'd247+xpc10nz) || (6'd61/*MS*/==-9'd246+xpc10nz) || (6'd61/*MS*/==-9'd245
              +xpc10nz) || (6'd61/*MS*/==-9'd244+xpc10nz) || (6'd61/*MS*/==-9'd242+xpc10nz) || (6'd61/*MS*/==-9'd241+xpc10nz) || (6'd61
              /*MS*/==-9'd239+xpc10nz) || (6'd61/*MS*/==-9'd238+xpc10nz) || (6'd61/*MS*/==-9'd236+xpc10nz) || (6'd61/*MS*/==-9'd171+xpc10nz
              ) || (6'd61/*MS*/==-8'd106+xpc10nz) || (6'd61/*MS*/==-8'd105+xpc10nz) || (6'd61/*MS*/==-8'd104+xpc10nz) || (6'd61/*MS*/==
              -8'd103+xpc10nz) || (6'd61/*MS*/==-8'd102+xpc10nz) || (6'd61/*MS*/==-8'd101+xpc10nz) || (6'd61/*MS*/==-8'd100+xpc10nz) || 
              (6'd61/*MS*/==-8'd99+xpc10nz) || (6'd61/*MS*/==-8'd98+xpc10nz) || (6'd61/*MS*/==-8'd97+xpc10nz) || (6'd61/*MS*/==-8'd96
              +xpc10nz) || (6'd61/*MS*/==-8'd95+xpc10nz) || (6'd61/*MS*/==-8'd94+xpc10nz) || (6'd61/*MS*/==-8'd93+xpc10nz) || (6'd61/*MS*/==
              -8'd92+xpc10nz) || (6'd61/*MS*/==-8'd91+xpc10nz) || (6'd61/*MS*/==-8'd90+xpc10nz) || (6'd61/*MS*/==-8'd89+xpc10nz) || (6'd61
              /*MS*/==-8'd88+xpc10nz) || (6'd61/*MS*/==-8'd87+xpc10nz) || (6'd61/*MS*/==-8'd86+xpc10nz) || (6'd61/*MS*/==-8'd85+xpc10nz
              ) || (6'd61/*MS*/==-8'd84+xpc10nz) || (6'd61/*MS*/==-8'd83+xpc10nz) || (6'd61/*MS*/==-8'd82+xpc10nz) || (6'd61/*MS*/==-8'd65
              +xpc10nz) || (6'd61/*MS*/==-8'd64+xpc10nz) || (6'd61/*MS*/==-7'd59+xpc10nz) || (6'd61/*MS*/==-7'd50+xpc10nz) || (6'd61/*MS*/==
              -7'd37+xpc10nz) || (6'd61/*MS*/==-6'd20+xpc10nz) || (6'd61/*MS*/==-6'd19+xpc10nz) || (6'd61/*MS*/==-6'd18+xpc10nz) || (6'd61
              /*MS*/==-6'd17+xpc10nz) || (6'd61/*MS*/==-6'd16+xpc10nz) || (6'd61/*MS*/==-5'd15+xpc10nz) || (6'd61/*MS*/==-5'd14+xpc10nz
              ) || (6'd61/*MS*/==-5'd13+xpc10nz) || (6'd61/*MS*/==-5'd12+xpc10nz) || (6'd61/*MS*/==-5'd11+xpc10nz) || (6'd61/*MS*/==-5'd10
              +xpc10nz) || (6'd61/*MS*/==-5'd9+xpc10nz) || (6'd61/*MS*/==-5'd8+xpc10nz) || (6'd61/*MS*/==-4'd7+xpc10nz) || (6'd61/*MS*/==
              -4'd6+xpc10nz) || (6'd61/*MS*/==-4'd5+xpc10nz) || (6'd61/*MS*/==-4'd4+xpc10nz) || (6'd61/*MS*/==-3'd3+xpc10nz) || (6'd61
              /*MS*/==-3'd2+xpc10nz) || (6'd61/*MS*/==-2'd1+xpc10nz) || (xpc10nz==6'd61/*US*/)) && !xpc10_clear && !xpc10_stall;

               xpc10_trk60 <= ((6'd60/*MS*/==-11'd609+xpc10nz) || (6'd60/*MS*/==-11'd599+xpc10nz) || (6'd60/*MS*/==-11'd588+xpc10nz) || 
              (6'd60/*MS*/==-11'd576+xpc10nz) || (6'd60/*MS*/==-11'd571+xpc10nz) || (6'd60/*MS*/==-11'd565+xpc10nz) || (6'd60/*MS*/==
              -11'd558+xpc10nz) || (6'd60/*MS*/==-11'd550+xpc10nz) || (6'd60/*MS*/==-11'd549+xpc10nz) || (6'd60/*MS*/==-11'd547+xpc10nz
              ) || (6'd60/*MS*/==-11'd544+xpc10nz) || (6'd60/*MS*/==-11'd540+xpc10nz) || (6'd60/*MS*/==-11'd539+xpc10nz) || (6'd60/*MS*/==
              -11'd537+xpc10nz) || (6'd60/*MS*/==-11'd534+xpc10nz) || (6'd60/*MS*/==-11'd532+xpc10nz) || (6'd60/*MS*/==-11'd528+xpc10nz
              ) || (6'd60/*MS*/==-10'd503+xpc10nz) || (6'd60/*MS*/==-10'd502+xpc10nz) || (6'd60/*MS*/==-10'd472+xpc10nz) || (6'd60/*MS*/==
              -10'd407+xpc10nz) || (6'd60/*MS*/==-10'd342+xpc10nz) || (6'd60/*MS*/==-10'd341+xpc10nz) || (6'd60/*MS*/==-10'd340+xpc10nz
              ) || (6'd60/*MS*/==-10'd338+xpc10nz) || (6'd60/*MS*/==-10'd335+xpc10nz) || (6'd60/*MS*/==-10'd334+xpc10nz) || (6'd60/*MS*/==
              -10'd330+xpc10nz) || (6'd60/*MS*/==-10'd329+xpc10nz) || (6'd60/*MS*/==-10'd327+xpc10nz) || (6'd60/*MS*/==-10'd324+xpc10nz
              ) || (6'd60/*MS*/==-10'd323+xpc10nz) || (6'd60/*MS*/==-10'd322+xpc10nz) || (6'd60/*MS*/==-10'd321+xpc10nz) || (6'd60/*MS*/==
              -10'd320+xpc10nz) || (6'd60/*MS*/==-10'd319+xpc10nz) || (6'd60/*MS*/==-10'd318+xpc10nz) || (6'd60/*MS*/==-10'd314+xpc10nz
              ) || (6'd60/*MS*/==-10'd289+xpc10nz) || (6'd60/*MS*/==-10'd287+xpc10nz) || (6'd60/*MS*/==-10'd285+xpc10nz) || (6'd60/*MS*/==
              -10'd284+xpc10nz) || (6'd60/*MS*/==-10'd259+xpc10nz) || (6'd60/*MS*/==-10'd258+xpc10nz) || (6'd60/*MS*/==-10'd257+xpc10nz
              ) || (6'd60/*MS*/==-9'd255+xpc10nz) || (6'd60/*MS*/==-9'd254+xpc10nz) || (6'd60/*MS*/==-9'd253+xpc10nz) || (6'd60/*MS*/==
              -9'd252+xpc10nz) || (6'd60/*MS*/==-9'd251+xpc10nz) || (6'd60/*MS*/==-9'd250+xpc10nz) || (6'd60/*MS*/==-9'd249+xpc10nz) || 
              (6'd60/*MS*/==-9'd248+xpc10nz) || (6'd60/*MS*/==-9'd247+xpc10nz) || (6'd60/*MS*/==-9'd246+xpc10nz) || (6'd60/*MS*/==-9'd245
              +xpc10nz) || (6'd60/*MS*/==-9'd244+xpc10nz) || (6'd60/*MS*/==-9'd242+xpc10nz) || (6'd60/*MS*/==-9'd241+xpc10nz) || (6'd60
              /*MS*/==-9'd239+xpc10nz) || (6'd60/*MS*/==-9'd238+xpc10nz) || (6'd60/*MS*/==-9'd236+xpc10nz) || (6'd60/*MS*/==-9'd171+xpc10nz
              ) || (6'd60/*MS*/==-8'd106+xpc10nz) || (6'd60/*MS*/==-8'd105+xpc10nz) || (6'd60/*MS*/==-8'd104+xpc10nz) || (6'd60/*MS*/==
              -8'd103+xpc10nz) || (6'd60/*MS*/==-8'd102+xpc10nz) || (6'd60/*MS*/==-8'd101+xpc10nz) || (6'd60/*MS*/==-8'd100+xpc10nz) || 
              (6'd60/*MS*/==-8'd99+xpc10nz) || (6'd60/*MS*/==-8'd98+xpc10nz) || (6'd60/*MS*/==-8'd97+xpc10nz) || (6'd60/*MS*/==-8'd96
              +xpc10nz) || (6'd60/*MS*/==-8'd95+xpc10nz) || (6'd60/*MS*/==-8'd94+xpc10nz) || (6'd60/*MS*/==-8'd93+xpc10nz) || (6'd60/*MS*/==
              -8'd92+xpc10nz) || (6'd60/*MS*/==-8'd91+xpc10nz) || (6'd60/*MS*/==-8'd90+xpc10nz) || (6'd60/*MS*/==-8'd89+xpc10nz) || (6'd60
              /*MS*/==-8'd88+xpc10nz) || (6'd60/*MS*/==-8'd87+xpc10nz) || (6'd60/*MS*/==-8'd86+xpc10nz) || (6'd60/*MS*/==-8'd85+xpc10nz
              ) || (6'd60/*MS*/==-8'd84+xpc10nz) || (6'd60/*MS*/==-8'd83+xpc10nz) || (6'd60/*MS*/==-8'd82+xpc10nz) || (6'd60/*MS*/==-8'd65
              +xpc10nz) || (6'd60/*MS*/==-8'd64+xpc10nz) || (6'd60/*MS*/==-7'd59+xpc10nz) || (6'd60/*MS*/==-7'd50+xpc10nz) || (6'd60/*MS*/==
              -7'd37+xpc10nz) || (6'd60/*MS*/==-6'd20+xpc10nz) || (6'd60/*MS*/==-6'd19+xpc10nz) || (6'd60/*MS*/==-6'd18+xpc10nz) || (6'd60
              /*MS*/==-6'd17+xpc10nz) || (6'd60/*MS*/==-6'd16+xpc10nz) || (6'd60/*MS*/==-5'd15+xpc10nz) || (6'd60/*MS*/==-5'd14+xpc10nz
              ) || (6'd60/*MS*/==-5'd13+xpc10nz) || (6'd60/*MS*/==-5'd12+xpc10nz) || (6'd60/*MS*/==-5'd11+xpc10nz) || (6'd60/*MS*/==-5'd10
              +xpc10nz) || (6'd60/*MS*/==-5'd9+xpc10nz) || (6'd60/*MS*/==-5'd8+xpc10nz) || (6'd60/*MS*/==-4'd7+xpc10nz) || (6'd60/*MS*/==
              -4'd6+xpc10nz) || (6'd60/*MS*/==-4'd5+xpc10nz) || (6'd60/*MS*/==-4'd4+xpc10nz) || (6'd60/*MS*/==-3'd3+xpc10nz) || (6'd60
              /*MS*/==-3'd2+xpc10nz) || (6'd60/*MS*/==-2'd1+xpc10nz) || (xpc10nz==6'd60/*US*/)) && !xpc10_clear && !xpc10_stall;

               xpc10_trk59 <= ((6'd59/*MS*/==-11'd609+xpc10nz) || (6'd59/*MS*/==-11'd599+xpc10nz) || (6'd59/*MS*/==-11'd588+xpc10nz) || 
              (6'd59/*MS*/==-11'd576+xpc10nz) || (6'd59/*MS*/==-11'd571+xpc10nz) || (6'd59/*MS*/==-11'd565+xpc10nz) || (6'd59/*MS*/==
              -11'd558+xpc10nz) || (6'd59/*MS*/==-11'd550+xpc10nz) || (6'd59/*MS*/==-11'd549+xpc10nz) || (6'd59/*MS*/==-11'd547+xpc10nz
              ) || (6'd59/*MS*/==-11'd544+xpc10nz) || (6'd59/*MS*/==-11'd540+xpc10nz) || (6'd59/*MS*/==-11'd539+xpc10nz) || (6'd59/*MS*/==
              -11'd537+xpc10nz) || (6'd59/*MS*/==-11'd534+xpc10nz) || (6'd59/*MS*/==-11'd532+xpc10nz) || (6'd59/*MS*/==-11'd528+xpc10nz
              ) || (6'd59/*MS*/==-10'd503+xpc10nz) || (6'd59/*MS*/==-10'd502+xpc10nz) || (6'd59/*MS*/==-10'd472+xpc10nz) || (6'd59/*MS*/==
              -10'd407+xpc10nz) || (6'd59/*MS*/==-10'd342+xpc10nz) || (6'd59/*MS*/==-10'd341+xpc10nz) || (6'd59/*MS*/==-10'd340+xpc10nz
              ) || (6'd59/*MS*/==-10'd338+xpc10nz) || (6'd59/*MS*/==-10'd335+xpc10nz) || (6'd59/*MS*/==-10'd334+xpc10nz) || (6'd59/*MS*/==
              -10'd330+xpc10nz) || (6'd59/*MS*/==-10'd329+xpc10nz) || (6'd59/*MS*/==-10'd327+xpc10nz) || (6'd59/*MS*/==-10'd324+xpc10nz
              ) || (6'd59/*MS*/==-10'd323+xpc10nz) || (6'd59/*MS*/==-10'd322+xpc10nz) || (6'd59/*MS*/==-10'd321+xpc10nz) || (6'd59/*MS*/==
              -10'd320+xpc10nz) || (6'd59/*MS*/==-10'd319+xpc10nz) || (6'd59/*MS*/==-10'd318+xpc10nz) || (6'd59/*MS*/==-10'd314+xpc10nz
              ) || (6'd59/*MS*/==-10'd289+xpc10nz) || (6'd59/*MS*/==-10'd287+xpc10nz) || (6'd59/*MS*/==-10'd285+xpc10nz) || (6'd59/*MS*/==
              -10'd284+xpc10nz) || (6'd59/*MS*/==-10'd259+xpc10nz) || (6'd59/*MS*/==-10'd258+xpc10nz) || (6'd59/*MS*/==-10'd257+xpc10nz
              ) || (6'd59/*MS*/==-9'd255+xpc10nz) || (6'd59/*MS*/==-9'd254+xpc10nz) || (6'd59/*MS*/==-9'd253+xpc10nz) || (6'd59/*MS*/==
              -9'd252+xpc10nz) || (6'd59/*MS*/==-9'd251+xpc10nz) || (6'd59/*MS*/==-9'd250+xpc10nz) || (6'd59/*MS*/==-9'd249+xpc10nz) || 
              (6'd59/*MS*/==-9'd248+xpc10nz) || (6'd59/*MS*/==-9'd247+xpc10nz) || (6'd59/*MS*/==-9'd246+xpc10nz) || (6'd59/*MS*/==-9'd245
              +xpc10nz) || (6'd59/*MS*/==-9'd244+xpc10nz) || (6'd59/*MS*/==-9'd242+xpc10nz) || (6'd59/*MS*/==-9'd241+xpc10nz) || (6'd59
              /*MS*/==-9'd239+xpc10nz) || (6'd59/*MS*/==-9'd238+xpc10nz) || (6'd59/*MS*/==-9'd236+xpc10nz) || (6'd59/*MS*/==-9'd171+xpc10nz
              ) || (6'd59/*MS*/==-8'd106+xpc10nz) || (6'd59/*MS*/==-8'd105+xpc10nz) || (6'd59/*MS*/==-8'd104+xpc10nz) || (6'd59/*MS*/==
              -8'd103+xpc10nz) || (6'd59/*MS*/==-8'd102+xpc10nz) || (6'd59/*MS*/==-8'd101+xpc10nz) || (6'd59/*MS*/==-8'd100+xpc10nz) || 
              (6'd59/*MS*/==-8'd99+xpc10nz) || (6'd59/*MS*/==-8'd98+xpc10nz) || (6'd59/*MS*/==-8'd97+xpc10nz) || (6'd59/*MS*/==-8'd96
              +xpc10nz) || (6'd59/*MS*/==-8'd95+xpc10nz) || (6'd59/*MS*/==-8'd94+xpc10nz) || (6'd59/*MS*/==-8'd93+xpc10nz) || (6'd59/*MS*/==
              -8'd92+xpc10nz) || (6'd59/*MS*/==-8'd91+xpc10nz) || (6'd59/*MS*/==-8'd90+xpc10nz) || (6'd59/*MS*/==-8'd89+xpc10nz) || (6'd59
              /*MS*/==-8'd88+xpc10nz) || (6'd59/*MS*/==-8'd87+xpc10nz) || (6'd59/*MS*/==-8'd86+xpc10nz) || (6'd59/*MS*/==-8'd85+xpc10nz
              ) || (6'd59/*MS*/==-8'd84+xpc10nz) || (6'd59/*MS*/==-8'd83+xpc10nz) || (6'd59/*MS*/==-8'd82+xpc10nz) || (6'd59/*MS*/==-8'd65
              +xpc10nz) || (6'd59/*MS*/==-8'd64+xpc10nz) || (6'd59/*MS*/==-7'd59+xpc10nz) || (6'd59/*MS*/==-7'd50+xpc10nz) || (6'd59/*MS*/==
              -7'd37+xpc10nz) || (6'd59/*MS*/==-6'd20+xpc10nz) || (6'd59/*MS*/==-6'd19+xpc10nz) || (6'd59/*MS*/==-6'd18+xpc10nz) || (6'd59
              /*MS*/==-6'd17+xpc10nz) || (6'd59/*MS*/==-6'd16+xpc10nz) || (6'd59/*MS*/==-5'd15+xpc10nz) || (6'd59/*MS*/==-5'd14+xpc10nz
              ) || (6'd59/*MS*/==-5'd13+xpc10nz) || (6'd59/*MS*/==-5'd12+xpc10nz) || (6'd59/*MS*/==-5'd11+xpc10nz) || (6'd59/*MS*/==-5'd10
              +xpc10nz) || (6'd59/*MS*/==-5'd9+xpc10nz) || (6'd59/*MS*/==-5'd8+xpc10nz) || (6'd59/*MS*/==-4'd7+xpc10nz) || (6'd59/*MS*/==
              -4'd6+xpc10nz) || (6'd59/*MS*/==-4'd5+xpc10nz) || (6'd59/*MS*/==-4'd4+xpc10nz) || (6'd59/*MS*/==-3'd3+xpc10nz) || (6'd59
              /*MS*/==-3'd2+xpc10nz) || (6'd59/*MS*/==-2'd1+xpc10nz) || (xpc10nz==6'd59/*US*/)) && !xpc10_clear && !xpc10_stall;

               xpc10_trk58 <= ((6'd58/*MS*/==-11'd609+xpc10nz) || (6'd58/*MS*/==-11'd599+xpc10nz) || (6'd58/*MS*/==-11'd588+xpc10nz) || 
              (6'd58/*MS*/==-11'd576+xpc10nz) || (6'd58/*MS*/==-11'd571+xpc10nz) || (6'd58/*MS*/==-11'd565+xpc10nz) || (6'd58/*MS*/==
              -11'd558+xpc10nz) || (6'd58/*MS*/==-11'd550+xpc10nz) || (6'd58/*MS*/==-11'd549+xpc10nz) || (6'd58/*MS*/==-11'd547+xpc10nz
              ) || (6'd58/*MS*/==-11'd544+xpc10nz) || (6'd58/*MS*/==-11'd540+xpc10nz) || (6'd58/*MS*/==-11'd539+xpc10nz) || (6'd58/*MS*/==
              -11'd537+xpc10nz) || (6'd58/*MS*/==-11'd534+xpc10nz) || (6'd58/*MS*/==-11'd532+xpc10nz) || (6'd58/*MS*/==-11'd528+xpc10nz
              ) || (6'd58/*MS*/==-10'd503+xpc10nz) || (6'd58/*MS*/==-10'd502+xpc10nz) || (6'd58/*MS*/==-10'd472+xpc10nz) || (6'd58/*MS*/==
              -10'd407+xpc10nz) || (6'd58/*MS*/==-10'd342+xpc10nz) || (6'd58/*MS*/==-10'd341+xpc10nz) || (6'd58/*MS*/==-10'd340+xpc10nz
              ) || (6'd58/*MS*/==-10'd338+xpc10nz) || (6'd58/*MS*/==-10'd335+xpc10nz) || (6'd58/*MS*/==-10'd334+xpc10nz) || (6'd58/*MS*/==
              -10'd330+xpc10nz) || (6'd58/*MS*/==-10'd329+xpc10nz) || (6'd58/*MS*/==-10'd327+xpc10nz) || (6'd58/*MS*/==-10'd324+xpc10nz
              ) || (6'd58/*MS*/==-10'd323+xpc10nz) || (6'd58/*MS*/==-10'd322+xpc10nz) || (6'd58/*MS*/==-10'd321+xpc10nz) || (6'd58/*MS*/==
              -10'd320+xpc10nz) || (6'd58/*MS*/==-10'd319+xpc10nz) || (6'd58/*MS*/==-10'd318+xpc10nz) || (6'd58/*MS*/==-10'd314+xpc10nz
              ) || (6'd58/*MS*/==-10'd289+xpc10nz) || (6'd58/*MS*/==-10'd287+xpc10nz) || (6'd58/*MS*/==-10'd285+xpc10nz) || (6'd58/*MS*/==
              -10'd284+xpc10nz) || (6'd58/*MS*/==-10'd259+xpc10nz) || (6'd58/*MS*/==-10'd258+xpc10nz) || (6'd58/*MS*/==-10'd257+xpc10nz
              ) || (6'd58/*MS*/==-9'd255+xpc10nz) || (6'd58/*MS*/==-9'd254+xpc10nz) || (6'd58/*MS*/==-9'd253+xpc10nz) || (6'd58/*MS*/==
              -9'd252+xpc10nz) || (6'd58/*MS*/==-9'd251+xpc10nz) || (6'd58/*MS*/==-9'd250+xpc10nz) || (6'd58/*MS*/==-9'd249+xpc10nz) || 
              (6'd58/*MS*/==-9'd248+xpc10nz) || (6'd58/*MS*/==-9'd247+xpc10nz) || (6'd58/*MS*/==-9'd246+xpc10nz) || (6'd58/*MS*/==-9'd245
              +xpc10nz) || (6'd58/*MS*/==-9'd244+xpc10nz) || (6'd58/*MS*/==-9'd242+xpc10nz) || (6'd58/*MS*/==-9'd241+xpc10nz) || (6'd58
              /*MS*/==-9'd239+xpc10nz) || (6'd58/*MS*/==-9'd238+xpc10nz) || (6'd58/*MS*/==-9'd236+xpc10nz) || (6'd58/*MS*/==-9'd171+xpc10nz
              ) || (6'd58/*MS*/==-8'd106+xpc10nz) || (6'd58/*MS*/==-8'd105+xpc10nz) || (6'd58/*MS*/==-8'd104+xpc10nz) || (6'd58/*MS*/==
              -8'd103+xpc10nz) || (6'd58/*MS*/==-8'd102+xpc10nz) || (6'd58/*MS*/==-8'd101+xpc10nz) || (6'd58/*MS*/==-8'd100+xpc10nz) || 
              (6'd58/*MS*/==-8'd99+xpc10nz) || (6'd58/*MS*/==-8'd98+xpc10nz) || (6'd58/*MS*/==-8'd97+xpc10nz) || (6'd58/*MS*/==-8'd96
              +xpc10nz) || (6'd58/*MS*/==-8'd95+xpc10nz) || (6'd58/*MS*/==-8'd94+xpc10nz) || (6'd58/*MS*/==-8'd93+xpc10nz) || (6'd58/*MS*/==
              -8'd92+xpc10nz) || (6'd58/*MS*/==-8'd91+xpc10nz) || (6'd58/*MS*/==-8'd90+xpc10nz) || (6'd58/*MS*/==-8'd89+xpc10nz) || (6'd58
              /*MS*/==-8'd88+xpc10nz) || (6'd58/*MS*/==-8'd87+xpc10nz) || (6'd58/*MS*/==-8'd86+xpc10nz) || (6'd58/*MS*/==-8'd85+xpc10nz
              ) || (6'd58/*MS*/==-8'd84+xpc10nz) || (6'd58/*MS*/==-8'd83+xpc10nz) || (6'd58/*MS*/==-8'd82+xpc10nz) || (6'd58/*MS*/==-8'd65
              +xpc10nz) || (6'd58/*MS*/==-8'd64+xpc10nz) || (6'd58/*MS*/==-7'd59+xpc10nz) || (6'd58/*MS*/==-7'd50+xpc10nz) || (6'd58/*MS*/==
              -7'd37+xpc10nz) || (6'd58/*MS*/==-6'd20+xpc10nz) || (6'd58/*MS*/==-6'd19+xpc10nz) || (6'd58/*MS*/==-6'd18+xpc10nz) || (6'd58
              /*MS*/==-6'd17+xpc10nz) || (6'd58/*MS*/==-6'd16+xpc10nz) || (6'd58/*MS*/==-5'd15+xpc10nz) || (6'd58/*MS*/==-5'd14+xpc10nz
              ) || (6'd58/*MS*/==-5'd13+xpc10nz) || (6'd58/*MS*/==-5'd12+xpc10nz) || (6'd58/*MS*/==-5'd11+xpc10nz) || (6'd58/*MS*/==-5'd10
              +xpc10nz) || (6'd58/*MS*/==-5'd9+xpc10nz) || (6'd58/*MS*/==-5'd8+xpc10nz) || (6'd58/*MS*/==-4'd7+xpc10nz) || (6'd58/*MS*/==
              -4'd6+xpc10nz) || (6'd58/*MS*/==-4'd5+xpc10nz) || (6'd58/*MS*/==-4'd4+xpc10nz) || (6'd58/*MS*/==-3'd3+xpc10nz) || (6'd58
              /*MS*/==-3'd2+xpc10nz) || (6'd58/*MS*/==-2'd1+xpc10nz) || (xpc10nz==6'd58/*US*/)) && !xpc10_clear && !xpc10_stall;

               xpc10_trk57 <= ((6'd57/*MS*/==-11'd609+xpc10nz) || (6'd57/*MS*/==-11'd599+xpc10nz) || (6'd57/*MS*/==-11'd588+xpc10nz) || 
              (6'd57/*MS*/==-11'd576+xpc10nz) || (6'd57/*MS*/==-11'd571+xpc10nz) || (6'd57/*MS*/==-11'd565+xpc10nz) || (6'd57/*MS*/==
              -11'd558+xpc10nz) || (6'd57/*MS*/==-11'd550+xpc10nz) || (6'd57/*MS*/==-11'd549+xpc10nz) || (6'd57/*MS*/==-11'd547+xpc10nz
              ) || (6'd57/*MS*/==-11'd544+xpc10nz) || (6'd57/*MS*/==-11'd540+xpc10nz) || (6'd57/*MS*/==-11'd539+xpc10nz) || (6'd57/*MS*/==
              -11'd537+xpc10nz) || (6'd57/*MS*/==-11'd534+xpc10nz) || (6'd57/*MS*/==-11'd532+xpc10nz) || (6'd57/*MS*/==-11'd528+xpc10nz
              ) || (6'd57/*MS*/==-10'd503+xpc10nz) || (6'd57/*MS*/==-10'd502+xpc10nz) || (6'd57/*MS*/==-10'd472+xpc10nz) || (6'd57/*MS*/==
              -10'd407+xpc10nz) || (6'd57/*MS*/==-10'd342+xpc10nz) || (6'd57/*MS*/==-10'd341+xpc10nz) || (6'd57/*MS*/==-10'd340+xpc10nz
              ) || (6'd57/*MS*/==-10'd338+xpc10nz) || (6'd57/*MS*/==-10'd335+xpc10nz) || (6'd57/*MS*/==-10'd334+xpc10nz) || (6'd57/*MS*/==
              -10'd330+xpc10nz) || (6'd57/*MS*/==-10'd329+xpc10nz) || (6'd57/*MS*/==-10'd327+xpc10nz) || (6'd57/*MS*/==-10'd324+xpc10nz
              ) || (6'd57/*MS*/==-10'd323+xpc10nz) || (6'd57/*MS*/==-10'd322+xpc10nz) || (6'd57/*MS*/==-10'd321+xpc10nz) || (6'd57/*MS*/==
              -10'd320+xpc10nz) || (6'd57/*MS*/==-10'd319+xpc10nz) || (6'd57/*MS*/==-10'd318+xpc10nz) || (6'd57/*MS*/==-10'd314+xpc10nz
              ) || (6'd57/*MS*/==-10'd289+xpc10nz) || (6'd57/*MS*/==-10'd287+xpc10nz) || (6'd57/*MS*/==-10'd285+xpc10nz) || (6'd57/*MS*/==
              -10'd284+xpc10nz) || (6'd57/*MS*/==-10'd259+xpc10nz) || (6'd57/*MS*/==-10'd258+xpc10nz) || (6'd57/*MS*/==-10'd257+xpc10nz
              ) || (6'd57/*MS*/==-9'd255+xpc10nz) || (6'd57/*MS*/==-9'd254+xpc10nz) || (6'd57/*MS*/==-9'd253+xpc10nz) || (6'd57/*MS*/==
              -9'd252+xpc10nz) || (6'd57/*MS*/==-9'd251+xpc10nz) || (6'd57/*MS*/==-9'd250+xpc10nz) || (6'd57/*MS*/==-9'd249+xpc10nz) || 
              (6'd57/*MS*/==-9'd248+xpc10nz) || (6'd57/*MS*/==-9'd247+xpc10nz) || (6'd57/*MS*/==-9'd246+xpc10nz) || (6'd57/*MS*/==-9'd245
              +xpc10nz) || (6'd57/*MS*/==-9'd244+xpc10nz) || (6'd57/*MS*/==-9'd242+xpc10nz) || (6'd57/*MS*/==-9'd241+xpc10nz) || (6'd57
              /*MS*/==-9'd239+xpc10nz) || (6'd57/*MS*/==-9'd238+xpc10nz) || (6'd57/*MS*/==-9'd236+xpc10nz) || (6'd57/*MS*/==-9'd171+xpc10nz
              ) || (6'd57/*MS*/==-8'd106+xpc10nz) || (6'd57/*MS*/==-8'd105+xpc10nz) || (6'd57/*MS*/==-8'd104+xpc10nz) || (6'd57/*MS*/==
              -8'd103+xpc10nz) || (6'd57/*MS*/==-8'd102+xpc10nz) || (6'd57/*MS*/==-8'd101+xpc10nz) || (6'd57/*MS*/==-8'd100+xpc10nz) || 
              (6'd57/*MS*/==-8'd99+xpc10nz) || (6'd57/*MS*/==-8'd98+xpc10nz) || (6'd57/*MS*/==-8'd97+xpc10nz) || (6'd57/*MS*/==-8'd96
              +xpc10nz) || (6'd57/*MS*/==-8'd95+xpc10nz) || (6'd57/*MS*/==-8'd94+xpc10nz) || (6'd57/*MS*/==-8'd93+xpc10nz) || (6'd57/*MS*/==
              -8'd92+xpc10nz) || (6'd57/*MS*/==-8'd91+xpc10nz) || (6'd57/*MS*/==-8'd90+xpc10nz) || (6'd57/*MS*/==-8'd89+xpc10nz) || (6'd57
              /*MS*/==-8'd88+xpc10nz) || (6'd57/*MS*/==-8'd87+xpc10nz) || (6'd57/*MS*/==-8'd86+xpc10nz) || (6'd57/*MS*/==-8'd85+xpc10nz
              ) || (6'd57/*MS*/==-8'd84+xpc10nz) || (6'd57/*MS*/==-8'd83+xpc10nz) || (6'd57/*MS*/==-8'd82+xpc10nz) || (6'd57/*MS*/==-8'd65
              +xpc10nz) || (6'd57/*MS*/==-8'd64+xpc10nz) || (6'd57/*MS*/==-7'd59+xpc10nz) || (6'd57/*MS*/==-7'd50+xpc10nz) || (6'd57/*MS*/==
              -7'd37+xpc10nz) || (6'd57/*MS*/==-6'd20+xpc10nz) || (6'd57/*MS*/==-6'd19+xpc10nz) || (6'd57/*MS*/==-6'd18+xpc10nz) || (6'd57
              /*MS*/==-6'd17+xpc10nz) || (6'd57/*MS*/==-6'd16+xpc10nz) || (6'd57/*MS*/==-5'd15+xpc10nz) || (6'd57/*MS*/==-5'd14+xpc10nz
              ) || (6'd57/*MS*/==-5'd13+xpc10nz) || (6'd57/*MS*/==-5'd12+xpc10nz) || (6'd57/*MS*/==-5'd11+xpc10nz) || (6'd57/*MS*/==-5'd10
              +xpc10nz) || (6'd57/*MS*/==-5'd9+xpc10nz) || (6'd57/*MS*/==-5'd8+xpc10nz) || (6'd57/*MS*/==-4'd7+xpc10nz) || (6'd57/*MS*/==
              -4'd6+xpc10nz) || (6'd57/*MS*/==-4'd5+xpc10nz) || (6'd57/*MS*/==-4'd4+xpc10nz) || (6'd57/*MS*/==-3'd3+xpc10nz) || (6'd57
              /*MS*/==-3'd2+xpc10nz) || (6'd57/*MS*/==-2'd1+xpc10nz) || (xpc10nz==6'd57/*US*/)) && !xpc10_clear && !xpc10_stall;

               xpc10_trk56 <= ((6'd56/*MS*/==-11'd609+xpc10nz) || (6'd56/*MS*/==-11'd599+xpc10nz) || (6'd56/*MS*/==-11'd588+xpc10nz) || 
              (6'd56/*MS*/==-11'd576+xpc10nz) || (6'd56/*MS*/==-11'd571+xpc10nz) || (6'd56/*MS*/==-11'd565+xpc10nz) || (6'd56/*MS*/==
              -11'd558+xpc10nz) || (6'd56/*MS*/==-11'd550+xpc10nz) || (6'd56/*MS*/==-11'd549+xpc10nz) || (6'd56/*MS*/==-11'd547+xpc10nz
              ) || (6'd56/*MS*/==-11'd544+xpc10nz) || (6'd56/*MS*/==-11'd540+xpc10nz) || (6'd56/*MS*/==-11'd539+xpc10nz) || (6'd56/*MS*/==
              -11'd537+xpc10nz) || (6'd56/*MS*/==-11'd534+xpc10nz) || (6'd56/*MS*/==-11'd532+xpc10nz) || (6'd56/*MS*/==-11'd528+xpc10nz
              ) || (6'd56/*MS*/==-10'd503+xpc10nz) || (6'd56/*MS*/==-10'd502+xpc10nz) || (6'd56/*MS*/==-10'd472+xpc10nz) || (6'd56/*MS*/==
              -10'd407+xpc10nz) || (6'd56/*MS*/==-10'd342+xpc10nz) || (6'd56/*MS*/==-10'd341+xpc10nz) || (6'd56/*MS*/==-10'd340+xpc10nz
              ) || (6'd56/*MS*/==-10'd338+xpc10nz) || (6'd56/*MS*/==-10'd335+xpc10nz) || (6'd56/*MS*/==-10'd334+xpc10nz) || (6'd56/*MS*/==
              -10'd330+xpc10nz) || (6'd56/*MS*/==-10'd329+xpc10nz) || (6'd56/*MS*/==-10'd327+xpc10nz) || (6'd56/*MS*/==-10'd324+xpc10nz
              ) || (6'd56/*MS*/==-10'd323+xpc10nz) || (6'd56/*MS*/==-10'd322+xpc10nz) || (6'd56/*MS*/==-10'd321+xpc10nz) || (6'd56/*MS*/==
              -10'd320+xpc10nz) || (6'd56/*MS*/==-10'd319+xpc10nz) || (6'd56/*MS*/==-10'd318+xpc10nz) || (6'd56/*MS*/==-10'd314+xpc10nz
              ) || (6'd56/*MS*/==-10'd289+xpc10nz) || (6'd56/*MS*/==-10'd287+xpc10nz) || (6'd56/*MS*/==-10'd285+xpc10nz) || (6'd56/*MS*/==
              -10'd284+xpc10nz) || (6'd56/*MS*/==-10'd259+xpc10nz) || (6'd56/*MS*/==-10'd258+xpc10nz) || (6'd56/*MS*/==-10'd257+xpc10nz
              ) || (6'd56/*MS*/==-9'd255+xpc10nz) || (6'd56/*MS*/==-9'd254+xpc10nz) || (6'd56/*MS*/==-9'd253+xpc10nz) || (6'd56/*MS*/==
              -9'd252+xpc10nz) || (6'd56/*MS*/==-9'd251+xpc10nz) || (6'd56/*MS*/==-9'd250+xpc10nz) || (6'd56/*MS*/==-9'd249+xpc10nz) || 
              (6'd56/*MS*/==-9'd248+xpc10nz) || (6'd56/*MS*/==-9'd247+xpc10nz) || (6'd56/*MS*/==-9'd246+xpc10nz) || (6'd56/*MS*/==-9'd245
              +xpc10nz) || (6'd56/*MS*/==-9'd244+xpc10nz) || (6'd56/*MS*/==-9'd242+xpc10nz) || (6'd56/*MS*/==-9'd241+xpc10nz) || (6'd56
              /*MS*/==-9'd239+xpc10nz) || (6'd56/*MS*/==-9'd238+xpc10nz) || (6'd56/*MS*/==-9'd236+xpc10nz) || (6'd56/*MS*/==-9'd171+xpc10nz
              ) || (6'd56/*MS*/==-8'd106+xpc10nz) || (6'd56/*MS*/==-8'd105+xpc10nz) || (6'd56/*MS*/==-8'd104+xpc10nz) || (6'd56/*MS*/==
              -8'd103+xpc10nz) || (6'd56/*MS*/==-8'd102+xpc10nz) || (6'd56/*MS*/==-8'd101+xpc10nz) || (6'd56/*MS*/==-8'd100+xpc10nz) || 
              (6'd56/*MS*/==-8'd99+xpc10nz) || (6'd56/*MS*/==-8'd98+xpc10nz) || (6'd56/*MS*/==-8'd97+xpc10nz) || (6'd56/*MS*/==-8'd96
              +xpc10nz) || (6'd56/*MS*/==-8'd95+xpc10nz) || (6'd56/*MS*/==-8'd94+xpc10nz) || (6'd56/*MS*/==-8'd93+xpc10nz) || (6'd56/*MS*/==
              -8'd92+xpc10nz) || (6'd56/*MS*/==-8'd91+xpc10nz) || (6'd56/*MS*/==-8'd90+xpc10nz) || (6'd56/*MS*/==-8'd89+xpc10nz) || (6'd56
              /*MS*/==-8'd88+xpc10nz) || (6'd56/*MS*/==-8'd87+xpc10nz) || (6'd56/*MS*/==-8'd86+xpc10nz) || (6'd56/*MS*/==-8'd85+xpc10nz
              ) || (6'd56/*MS*/==-8'd84+xpc10nz) || (6'd56/*MS*/==-8'd83+xpc10nz) || (6'd56/*MS*/==-8'd82+xpc10nz) || (6'd56/*MS*/==-8'd65
              +xpc10nz) || (6'd56/*MS*/==-8'd64+xpc10nz) || (6'd56/*MS*/==-7'd59+xpc10nz) || (6'd56/*MS*/==-7'd50+xpc10nz) || (6'd56/*MS*/==
              -7'd37+xpc10nz) || (6'd56/*MS*/==-6'd20+xpc10nz) || (6'd56/*MS*/==-6'd19+xpc10nz) || (6'd56/*MS*/==-6'd18+xpc10nz) || (6'd56
              /*MS*/==-6'd17+xpc10nz) || (6'd56/*MS*/==-6'd16+xpc10nz) || (6'd56/*MS*/==-5'd15+xpc10nz) || (6'd56/*MS*/==-5'd14+xpc10nz
              ) || (6'd56/*MS*/==-5'd13+xpc10nz) || (6'd56/*MS*/==-5'd12+xpc10nz) || (6'd56/*MS*/==-5'd11+xpc10nz) || (6'd56/*MS*/==-5'd10
              +xpc10nz) || (6'd56/*MS*/==-5'd9+xpc10nz) || (6'd56/*MS*/==-5'd8+xpc10nz) || (6'd56/*MS*/==-4'd7+xpc10nz) || (6'd56/*MS*/==
              -4'd6+xpc10nz) || (6'd56/*MS*/==-4'd5+xpc10nz) || (6'd56/*MS*/==-4'd4+xpc10nz) || (6'd56/*MS*/==-3'd3+xpc10nz) || (6'd56
              /*MS*/==-3'd2+xpc10nz) || (6'd56/*MS*/==-2'd1+xpc10nz) || (xpc10nz==6'd56/*US*/)) && !xpc10_clear && !xpc10_stall;

               xpc10_trk55 <= ((6'd55/*MS*/==-11'd609+xpc10nz) || (6'd55/*MS*/==-11'd599+xpc10nz) || (6'd55/*MS*/==-11'd588+xpc10nz) || 
              (6'd55/*MS*/==-11'd576+xpc10nz) || (6'd55/*MS*/==-11'd571+xpc10nz) || (6'd55/*MS*/==-11'd565+xpc10nz) || (6'd55/*MS*/==
              -11'd558+xpc10nz) || (6'd55/*MS*/==-11'd550+xpc10nz) || (6'd55/*MS*/==-11'd549+xpc10nz) || (6'd55/*MS*/==-11'd547+xpc10nz
              ) || (6'd55/*MS*/==-11'd544+xpc10nz) || (6'd55/*MS*/==-11'd540+xpc10nz) || (6'd55/*MS*/==-11'd539+xpc10nz) || (6'd55/*MS*/==
              -11'd537+xpc10nz) || (6'd55/*MS*/==-11'd534+xpc10nz) || (6'd55/*MS*/==-11'd532+xpc10nz) || (6'd55/*MS*/==-11'd528+xpc10nz
              ) || (6'd55/*MS*/==-10'd503+xpc10nz) || (6'd55/*MS*/==-10'd502+xpc10nz) || (6'd55/*MS*/==-10'd472+xpc10nz) || (6'd55/*MS*/==
              -10'd407+xpc10nz) || (6'd55/*MS*/==-10'd342+xpc10nz) || (6'd55/*MS*/==-10'd341+xpc10nz) || (6'd55/*MS*/==-10'd340+xpc10nz
              ) || (6'd55/*MS*/==-10'd338+xpc10nz) || (6'd55/*MS*/==-10'd335+xpc10nz) || (6'd55/*MS*/==-10'd334+xpc10nz) || (6'd55/*MS*/==
              -10'd330+xpc10nz) || (6'd55/*MS*/==-10'd329+xpc10nz) || (6'd55/*MS*/==-10'd327+xpc10nz) || (6'd55/*MS*/==-10'd324+xpc10nz
              ) || (6'd55/*MS*/==-10'd323+xpc10nz) || (6'd55/*MS*/==-10'd322+xpc10nz) || (6'd55/*MS*/==-10'd321+xpc10nz) || (6'd55/*MS*/==
              -10'd320+xpc10nz) || (6'd55/*MS*/==-10'd319+xpc10nz) || (6'd55/*MS*/==-10'd318+xpc10nz) || (6'd55/*MS*/==-10'd314+xpc10nz
              ) || (6'd55/*MS*/==-10'd289+xpc10nz) || (6'd55/*MS*/==-10'd287+xpc10nz) || (6'd55/*MS*/==-10'd285+xpc10nz) || (6'd55/*MS*/==
              -10'd284+xpc10nz) || (6'd55/*MS*/==-10'd259+xpc10nz) || (6'd55/*MS*/==-10'd258+xpc10nz) || (6'd55/*MS*/==-10'd257+xpc10nz
              ) || (6'd55/*MS*/==-9'd255+xpc10nz) || (6'd55/*MS*/==-9'd254+xpc10nz) || (6'd55/*MS*/==-9'd253+xpc10nz) || (6'd55/*MS*/==
              -9'd252+xpc10nz) || (6'd55/*MS*/==-9'd251+xpc10nz) || (6'd55/*MS*/==-9'd250+xpc10nz) || (6'd55/*MS*/==-9'd249+xpc10nz) || 
              (6'd55/*MS*/==-9'd248+xpc10nz) || (6'd55/*MS*/==-9'd247+xpc10nz) || (6'd55/*MS*/==-9'd246+xpc10nz) || (6'd55/*MS*/==-9'd245
              +xpc10nz) || (6'd55/*MS*/==-9'd244+xpc10nz) || (6'd55/*MS*/==-9'd242+xpc10nz) || (6'd55/*MS*/==-9'd241+xpc10nz) || (6'd55
              /*MS*/==-9'd239+xpc10nz) || (6'd55/*MS*/==-9'd238+xpc10nz) || (6'd55/*MS*/==-9'd236+xpc10nz) || (6'd55/*MS*/==-9'd171+xpc10nz
              ) || (6'd55/*MS*/==-8'd106+xpc10nz) || (6'd55/*MS*/==-8'd105+xpc10nz) || (6'd55/*MS*/==-8'd104+xpc10nz) || (6'd55/*MS*/==
              -8'd103+xpc10nz) || (6'd55/*MS*/==-8'd102+xpc10nz) || (6'd55/*MS*/==-8'd101+xpc10nz) || (6'd55/*MS*/==-8'd100+xpc10nz) || 
              (6'd55/*MS*/==-8'd99+xpc10nz) || (6'd55/*MS*/==-8'd98+xpc10nz) || (6'd55/*MS*/==-8'd97+xpc10nz) || (6'd55/*MS*/==-8'd96
              +xpc10nz) || (6'd55/*MS*/==-8'd95+xpc10nz) || (6'd55/*MS*/==-8'd94+xpc10nz) || (6'd55/*MS*/==-8'd93+xpc10nz) || (6'd55/*MS*/==
              -8'd92+xpc10nz) || (6'd55/*MS*/==-8'd91+xpc10nz) || (6'd55/*MS*/==-8'd90+xpc10nz) || (6'd55/*MS*/==-8'd89+xpc10nz) || (6'd55
              /*MS*/==-8'd88+xpc10nz) || (6'd55/*MS*/==-8'd87+xpc10nz) || (6'd55/*MS*/==-8'd86+xpc10nz) || (6'd55/*MS*/==-8'd85+xpc10nz
              ) || (6'd55/*MS*/==-8'd84+xpc10nz) || (6'd55/*MS*/==-8'd83+xpc10nz) || (6'd55/*MS*/==-8'd82+xpc10nz) || (6'd55/*MS*/==-8'd65
              +xpc10nz) || (6'd55/*MS*/==-8'd64+xpc10nz) || (6'd55/*MS*/==-7'd59+xpc10nz) || (6'd55/*MS*/==-7'd50+xpc10nz) || (6'd55/*MS*/==
              -7'd37+xpc10nz) || (6'd55/*MS*/==-6'd20+xpc10nz) || (6'd55/*MS*/==-6'd19+xpc10nz) || (6'd55/*MS*/==-6'd18+xpc10nz) || (6'd55
              /*MS*/==-6'd17+xpc10nz) || (6'd55/*MS*/==-6'd16+xpc10nz) || (6'd55/*MS*/==-5'd15+xpc10nz) || (6'd55/*MS*/==-5'd14+xpc10nz
              ) || (6'd55/*MS*/==-5'd13+xpc10nz) || (6'd55/*MS*/==-5'd12+xpc10nz) || (6'd55/*MS*/==-5'd11+xpc10nz) || (6'd55/*MS*/==-5'd10
              +xpc10nz) || (6'd55/*MS*/==-5'd9+xpc10nz) || (6'd55/*MS*/==-5'd8+xpc10nz) || (6'd55/*MS*/==-4'd7+xpc10nz) || (6'd55/*MS*/==
              -4'd6+xpc10nz) || (6'd55/*MS*/==-4'd5+xpc10nz) || (6'd55/*MS*/==-4'd4+xpc10nz) || (6'd55/*MS*/==-3'd3+xpc10nz) || (6'd55
              /*MS*/==-3'd2+xpc10nz) || (6'd55/*MS*/==-2'd1+xpc10nz) || (xpc10nz==6'd55/*US*/)) && !xpc10_clear && !xpc10_stall;

               xpc10_trk54 <= ((6'd54/*MS*/==-11'd609+xpc10nz) || (6'd54/*MS*/==-11'd599+xpc10nz) || (6'd54/*MS*/==-11'd588+xpc10nz) || 
              (6'd54/*MS*/==-11'd576+xpc10nz) || (6'd54/*MS*/==-11'd571+xpc10nz) || (6'd54/*MS*/==-11'd565+xpc10nz) || (6'd54/*MS*/==
              -11'd558+xpc10nz) || (6'd54/*MS*/==-11'd550+xpc10nz) || (6'd54/*MS*/==-11'd549+xpc10nz) || (6'd54/*MS*/==-11'd547+xpc10nz
              ) || (6'd54/*MS*/==-11'd544+xpc10nz) || (6'd54/*MS*/==-11'd540+xpc10nz) || (6'd54/*MS*/==-11'd539+xpc10nz) || (6'd54/*MS*/==
              -11'd537+xpc10nz) || (6'd54/*MS*/==-11'd534+xpc10nz) || (6'd54/*MS*/==-11'd532+xpc10nz) || (6'd54/*MS*/==-11'd528+xpc10nz
              ) || (6'd54/*MS*/==-10'd503+xpc10nz) || (6'd54/*MS*/==-10'd502+xpc10nz) || (6'd54/*MS*/==-10'd472+xpc10nz) || (6'd54/*MS*/==
              -10'd407+xpc10nz) || (6'd54/*MS*/==-10'd342+xpc10nz) || (6'd54/*MS*/==-10'd341+xpc10nz) || (6'd54/*MS*/==-10'd340+xpc10nz
              ) || (6'd54/*MS*/==-10'd338+xpc10nz) || (6'd54/*MS*/==-10'd335+xpc10nz) || (6'd54/*MS*/==-10'd334+xpc10nz) || (6'd54/*MS*/==
              -10'd330+xpc10nz) || (6'd54/*MS*/==-10'd329+xpc10nz) || (6'd54/*MS*/==-10'd327+xpc10nz) || (6'd54/*MS*/==-10'd324+xpc10nz
              ) || (6'd54/*MS*/==-10'd323+xpc10nz) || (6'd54/*MS*/==-10'd322+xpc10nz) || (6'd54/*MS*/==-10'd321+xpc10nz) || (6'd54/*MS*/==
              -10'd320+xpc10nz) || (6'd54/*MS*/==-10'd319+xpc10nz) || (6'd54/*MS*/==-10'd318+xpc10nz) || (6'd54/*MS*/==-10'd314+xpc10nz
              ) || (6'd54/*MS*/==-10'd289+xpc10nz) || (6'd54/*MS*/==-10'd287+xpc10nz) || (6'd54/*MS*/==-10'd285+xpc10nz) || (6'd54/*MS*/==
              -10'd284+xpc10nz) || (6'd54/*MS*/==-10'd259+xpc10nz) || (6'd54/*MS*/==-10'd258+xpc10nz) || (6'd54/*MS*/==-10'd257+xpc10nz
              ) || (6'd54/*MS*/==-9'd255+xpc10nz) || (6'd54/*MS*/==-9'd254+xpc10nz) || (6'd54/*MS*/==-9'd253+xpc10nz) || (6'd54/*MS*/==
              -9'd252+xpc10nz) || (6'd54/*MS*/==-9'd251+xpc10nz) || (6'd54/*MS*/==-9'd250+xpc10nz) || (6'd54/*MS*/==-9'd249+xpc10nz) || 
              (6'd54/*MS*/==-9'd248+xpc10nz) || (6'd54/*MS*/==-9'd247+xpc10nz) || (6'd54/*MS*/==-9'd246+xpc10nz) || (6'd54/*MS*/==-9'd245
              +xpc10nz) || (6'd54/*MS*/==-9'd244+xpc10nz) || (6'd54/*MS*/==-9'd242+xpc10nz) || (6'd54/*MS*/==-9'd241+xpc10nz) || (6'd54
              /*MS*/==-9'd239+xpc10nz) || (6'd54/*MS*/==-9'd238+xpc10nz) || (6'd54/*MS*/==-9'd236+xpc10nz) || (6'd54/*MS*/==-9'd171+xpc10nz
              ) || (6'd54/*MS*/==-8'd106+xpc10nz) || (6'd54/*MS*/==-8'd105+xpc10nz) || (6'd54/*MS*/==-8'd104+xpc10nz) || (6'd54/*MS*/==
              -8'd103+xpc10nz) || (6'd54/*MS*/==-8'd102+xpc10nz) || (6'd54/*MS*/==-8'd101+xpc10nz) || (6'd54/*MS*/==-8'd100+xpc10nz) || 
              (6'd54/*MS*/==-8'd99+xpc10nz) || (6'd54/*MS*/==-8'd98+xpc10nz) || (6'd54/*MS*/==-8'd97+xpc10nz) || (6'd54/*MS*/==-8'd96
              +xpc10nz) || (6'd54/*MS*/==-8'd95+xpc10nz) || (6'd54/*MS*/==-8'd94+xpc10nz) || (6'd54/*MS*/==-8'd93+xpc10nz) || (6'd54/*MS*/==
              -8'd92+xpc10nz) || (6'd54/*MS*/==-8'd91+xpc10nz) || (6'd54/*MS*/==-8'd90+xpc10nz) || (6'd54/*MS*/==-8'd89+xpc10nz) || (6'd54
              /*MS*/==-8'd88+xpc10nz) || (6'd54/*MS*/==-8'd87+xpc10nz) || (6'd54/*MS*/==-8'd86+xpc10nz) || (6'd54/*MS*/==-8'd85+xpc10nz
              ) || (6'd54/*MS*/==-8'd84+xpc10nz) || (6'd54/*MS*/==-8'd83+xpc10nz) || (6'd54/*MS*/==-8'd82+xpc10nz) || (6'd54/*MS*/==-8'd65
              +xpc10nz) || (6'd54/*MS*/==-8'd64+xpc10nz) || (6'd54/*MS*/==-7'd59+xpc10nz) || (6'd54/*MS*/==-7'd50+xpc10nz) || (6'd54/*MS*/==
              -7'd37+xpc10nz) || (6'd54/*MS*/==-6'd20+xpc10nz) || (6'd54/*MS*/==-6'd19+xpc10nz) || (6'd54/*MS*/==-6'd18+xpc10nz) || (6'd54
              /*MS*/==-6'd17+xpc10nz) || (6'd54/*MS*/==-6'd16+xpc10nz) || (6'd54/*MS*/==-5'd15+xpc10nz) || (6'd54/*MS*/==-5'd14+xpc10nz
              ) || (6'd54/*MS*/==-5'd13+xpc10nz) || (6'd54/*MS*/==-5'd12+xpc10nz) || (6'd54/*MS*/==-5'd11+xpc10nz) || (6'd54/*MS*/==-5'd10
              +xpc10nz) || (6'd54/*MS*/==-5'd9+xpc10nz) || (6'd54/*MS*/==-5'd8+xpc10nz) || (6'd54/*MS*/==-4'd7+xpc10nz) || (6'd54/*MS*/==
              -4'd6+xpc10nz) || (6'd54/*MS*/==-4'd5+xpc10nz) || (6'd54/*MS*/==-4'd4+xpc10nz) || (6'd54/*MS*/==-3'd3+xpc10nz) || (6'd54
              /*MS*/==-3'd2+xpc10nz) || (6'd54/*MS*/==-2'd1+xpc10nz) || (xpc10nz==6'd54/*US*/)) && !xpc10_clear && !xpc10_stall;

               xpc10_trk53 <= ((6'd53/*MS*/==-11'd609+xpc10nz) || (6'd53/*MS*/==-11'd599+xpc10nz) || (6'd53/*MS*/==-11'd588+xpc10nz) || 
              (6'd53/*MS*/==-11'd576+xpc10nz) || (6'd53/*MS*/==-11'd571+xpc10nz) || (6'd53/*MS*/==-11'd565+xpc10nz) || (6'd53/*MS*/==
              -11'd558+xpc10nz) || (6'd53/*MS*/==-11'd550+xpc10nz) || (6'd53/*MS*/==-11'd549+xpc10nz) || (6'd53/*MS*/==-11'd547+xpc10nz
              ) || (6'd53/*MS*/==-11'd544+xpc10nz) || (6'd53/*MS*/==-11'd540+xpc10nz) || (6'd53/*MS*/==-11'd539+xpc10nz) || (6'd53/*MS*/==
              -11'd537+xpc10nz) || (6'd53/*MS*/==-11'd534+xpc10nz) || (6'd53/*MS*/==-11'd532+xpc10nz) || (6'd53/*MS*/==-11'd528+xpc10nz
              ) || (6'd53/*MS*/==-10'd503+xpc10nz) || (6'd53/*MS*/==-10'd502+xpc10nz) || (6'd53/*MS*/==-10'd472+xpc10nz) || (6'd53/*MS*/==
              -10'd407+xpc10nz) || (6'd53/*MS*/==-10'd342+xpc10nz) || (6'd53/*MS*/==-10'd341+xpc10nz) || (6'd53/*MS*/==-10'd340+xpc10nz
              ) || (6'd53/*MS*/==-10'd338+xpc10nz) || (6'd53/*MS*/==-10'd335+xpc10nz) || (6'd53/*MS*/==-10'd334+xpc10nz) || (6'd53/*MS*/==
              -10'd330+xpc10nz) || (6'd53/*MS*/==-10'd329+xpc10nz) || (6'd53/*MS*/==-10'd327+xpc10nz) || (6'd53/*MS*/==-10'd324+xpc10nz
              ) || (6'd53/*MS*/==-10'd323+xpc10nz) || (6'd53/*MS*/==-10'd322+xpc10nz) || (6'd53/*MS*/==-10'd321+xpc10nz) || (6'd53/*MS*/==
              -10'd320+xpc10nz) || (6'd53/*MS*/==-10'd319+xpc10nz) || (6'd53/*MS*/==-10'd318+xpc10nz) || (6'd53/*MS*/==-10'd314+xpc10nz
              ) || (6'd53/*MS*/==-10'd289+xpc10nz) || (6'd53/*MS*/==-10'd287+xpc10nz) || (6'd53/*MS*/==-10'd285+xpc10nz) || (6'd53/*MS*/==
              -10'd284+xpc10nz) || (6'd53/*MS*/==-10'd259+xpc10nz) || (6'd53/*MS*/==-10'd258+xpc10nz) || (6'd53/*MS*/==-10'd257+xpc10nz
              ) || (6'd53/*MS*/==-9'd255+xpc10nz) || (6'd53/*MS*/==-9'd254+xpc10nz) || (6'd53/*MS*/==-9'd253+xpc10nz) || (6'd53/*MS*/==
              -9'd252+xpc10nz) || (6'd53/*MS*/==-9'd251+xpc10nz) || (6'd53/*MS*/==-9'd250+xpc10nz) || (6'd53/*MS*/==-9'd249+xpc10nz) || 
              (6'd53/*MS*/==-9'd248+xpc10nz) || (6'd53/*MS*/==-9'd247+xpc10nz) || (6'd53/*MS*/==-9'd246+xpc10nz) || (6'd53/*MS*/==-9'd245
              +xpc10nz) || (6'd53/*MS*/==-9'd244+xpc10nz) || (6'd53/*MS*/==-9'd242+xpc10nz) || (6'd53/*MS*/==-9'd241+xpc10nz) || (6'd53
              /*MS*/==-9'd239+xpc10nz) || (6'd53/*MS*/==-9'd238+xpc10nz) || (6'd53/*MS*/==-9'd236+xpc10nz) || (6'd53/*MS*/==-9'd171+xpc10nz
              ) || (6'd53/*MS*/==-8'd106+xpc10nz) || (6'd53/*MS*/==-8'd105+xpc10nz) || (6'd53/*MS*/==-8'd104+xpc10nz) || (6'd53/*MS*/==
              -8'd103+xpc10nz) || (6'd53/*MS*/==-8'd102+xpc10nz) || (6'd53/*MS*/==-8'd101+xpc10nz) || (6'd53/*MS*/==-8'd100+xpc10nz) || 
              (6'd53/*MS*/==-8'd99+xpc10nz) || (6'd53/*MS*/==-8'd98+xpc10nz) || (6'd53/*MS*/==-8'd97+xpc10nz) || (6'd53/*MS*/==-8'd96
              +xpc10nz) || (6'd53/*MS*/==-8'd95+xpc10nz) || (6'd53/*MS*/==-8'd94+xpc10nz) || (6'd53/*MS*/==-8'd93+xpc10nz) || (6'd53/*MS*/==
              -8'd92+xpc10nz) || (6'd53/*MS*/==-8'd91+xpc10nz) || (6'd53/*MS*/==-8'd90+xpc10nz) || (6'd53/*MS*/==-8'd89+xpc10nz) || (6'd53
              /*MS*/==-8'd88+xpc10nz) || (6'd53/*MS*/==-8'd87+xpc10nz) || (6'd53/*MS*/==-8'd86+xpc10nz) || (6'd53/*MS*/==-8'd85+xpc10nz
              ) || (6'd53/*MS*/==-8'd84+xpc10nz) || (6'd53/*MS*/==-8'd83+xpc10nz) || (6'd53/*MS*/==-8'd82+xpc10nz) || (6'd53/*MS*/==-8'd65
              +xpc10nz) || (6'd53/*MS*/==-8'd64+xpc10nz) || (6'd53/*MS*/==-7'd59+xpc10nz) || (6'd53/*MS*/==-7'd50+xpc10nz) || (6'd53/*MS*/==
              -7'd37+xpc10nz) || (6'd53/*MS*/==-6'd20+xpc10nz) || (6'd53/*MS*/==-6'd19+xpc10nz) || (6'd53/*MS*/==-6'd18+xpc10nz) || (6'd53
              /*MS*/==-6'd17+xpc10nz) || (6'd53/*MS*/==-6'd16+xpc10nz) || (6'd53/*MS*/==-5'd15+xpc10nz) || (6'd53/*MS*/==-5'd14+xpc10nz
              ) || (6'd53/*MS*/==-5'd13+xpc10nz) || (6'd53/*MS*/==-5'd12+xpc10nz) || (6'd53/*MS*/==-5'd11+xpc10nz) || (6'd53/*MS*/==-5'd10
              +xpc10nz) || (6'd53/*MS*/==-5'd9+xpc10nz) || (6'd53/*MS*/==-5'd8+xpc10nz) || (6'd53/*MS*/==-4'd7+xpc10nz) || (6'd53/*MS*/==
              -4'd6+xpc10nz) || (6'd53/*MS*/==-4'd5+xpc10nz) || (6'd53/*MS*/==-4'd4+xpc10nz) || (6'd53/*MS*/==-3'd3+xpc10nz) || (6'd53
              /*MS*/==-3'd2+xpc10nz) || (6'd53/*MS*/==-2'd1+xpc10nz) || (xpc10nz==6'd53/*US*/)) && !xpc10_clear && !xpc10_stall;

               xpc10_trk52 <= ((6'd52/*MS*/==-11'd609+xpc10nz) || (6'd52/*MS*/==-11'd599+xpc10nz) || (6'd52/*MS*/==-11'd588+xpc10nz) || 
              (6'd52/*MS*/==-11'd576+xpc10nz) || (6'd52/*MS*/==-11'd571+xpc10nz) || (6'd52/*MS*/==-11'd565+xpc10nz) || (6'd52/*MS*/==
              -11'd558+xpc10nz) || (6'd52/*MS*/==-11'd550+xpc10nz) || (6'd52/*MS*/==-11'd549+xpc10nz) || (6'd52/*MS*/==-11'd547+xpc10nz
              ) || (6'd52/*MS*/==-11'd544+xpc10nz) || (6'd52/*MS*/==-11'd540+xpc10nz) || (6'd52/*MS*/==-11'd539+xpc10nz) || (6'd52/*MS*/==
              -11'd537+xpc10nz) || (6'd52/*MS*/==-11'd534+xpc10nz) || (6'd52/*MS*/==-11'd532+xpc10nz) || (6'd52/*MS*/==-11'd528+xpc10nz
              ) || (6'd52/*MS*/==-10'd503+xpc10nz) || (6'd52/*MS*/==-10'd502+xpc10nz) || (6'd52/*MS*/==-10'd472+xpc10nz) || (6'd52/*MS*/==
              -10'd407+xpc10nz) || (6'd52/*MS*/==-10'd342+xpc10nz) || (6'd52/*MS*/==-10'd341+xpc10nz) || (6'd52/*MS*/==-10'd340+xpc10nz
              ) || (6'd52/*MS*/==-10'd338+xpc10nz) || (6'd52/*MS*/==-10'd335+xpc10nz) || (6'd52/*MS*/==-10'd334+xpc10nz) || (6'd52/*MS*/==
              -10'd330+xpc10nz) || (6'd52/*MS*/==-10'd329+xpc10nz) || (6'd52/*MS*/==-10'd327+xpc10nz) || (6'd52/*MS*/==-10'd324+xpc10nz
              ) || (6'd52/*MS*/==-10'd323+xpc10nz) || (6'd52/*MS*/==-10'd322+xpc10nz) || (6'd52/*MS*/==-10'd321+xpc10nz) || (6'd52/*MS*/==
              -10'd320+xpc10nz) || (6'd52/*MS*/==-10'd319+xpc10nz) || (6'd52/*MS*/==-10'd318+xpc10nz) || (6'd52/*MS*/==-10'd314+xpc10nz
              ) || (6'd52/*MS*/==-10'd289+xpc10nz) || (6'd52/*MS*/==-10'd287+xpc10nz) || (6'd52/*MS*/==-10'd285+xpc10nz) || (6'd52/*MS*/==
              -10'd284+xpc10nz) || (6'd52/*MS*/==-10'd259+xpc10nz) || (6'd52/*MS*/==-10'd258+xpc10nz) || (6'd52/*MS*/==-10'd257+xpc10nz
              ) || (6'd52/*MS*/==-9'd255+xpc10nz) || (6'd52/*MS*/==-9'd254+xpc10nz) || (6'd52/*MS*/==-9'd253+xpc10nz) || (6'd52/*MS*/==
              -9'd252+xpc10nz) || (6'd52/*MS*/==-9'd251+xpc10nz) || (6'd52/*MS*/==-9'd250+xpc10nz) || (6'd52/*MS*/==-9'd249+xpc10nz) || 
              (6'd52/*MS*/==-9'd248+xpc10nz) || (6'd52/*MS*/==-9'd247+xpc10nz) || (6'd52/*MS*/==-9'd246+xpc10nz) || (6'd52/*MS*/==-9'd245
              +xpc10nz) || (6'd52/*MS*/==-9'd244+xpc10nz) || (6'd52/*MS*/==-9'd242+xpc10nz) || (6'd52/*MS*/==-9'd241+xpc10nz) || (6'd52
              /*MS*/==-9'd239+xpc10nz) || (6'd52/*MS*/==-9'd238+xpc10nz) || (6'd52/*MS*/==-9'd236+xpc10nz) || (6'd52/*MS*/==-9'd171+xpc10nz
              ) || (6'd52/*MS*/==-8'd106+xpc10nz) || (6'd52/*MS*/==-8'd105+xpc10nz) || (6'd52/*MS*/==-8'd104+xpc10nz) || (6'd52/*MS*/==
              -8'd103+xpc10nz) || (6'd52/*MS*/==-8'd102+xpc10nz) || (6'd52/*MS*/==-8'd101+xpc10nz) || (6'd52/*MS*/==-8'd100+xpc10nz) || 
              (6'd52/*MS*/==-8'd99+xpc10nz) || (6'd52/*MS*/==-8'd98+xpc10nz) || (6'd52/*MS*/==-8'd97+xpc10nz) || (6'd52/*MS*/==-8'd96
              +xpc10nz) || (6'd52/*MS*/==-8'd95+xpc10nz) || (6'd52/*MS*/==-8'd94+xpc10nz) || (6'd52/*MS*/==-8'd93+xpc10nz) || (6'd52/*MS*/==
              -8'd92+xpc10nz) || (6'd52/*MS*/==-8'd91+xpc10nz) || (6'd52/*MS*/==-8'd90+xpc10nz) || (6'd52/*MS*/==-8'd89+xpc10nz) || (6'd52
              /*MS*/==-8'd88+xpc10nz) || (6'd52/*MS*/==-8'd87+xpc10nz) || (6'd52/*MS*/==-8'd86+xpc10nz) || (6'd52/*MS*/==-8'd85+xpc10nz
              ) || (6'd52/*MS*/==-8'd84+xpc10nz) || (6'd52/*MS*/==-8'd83+xpc10nz) || (6'd52/*MS*/==-8'd82+xpc10nz) || (6'd52/*MS*/==-8'd65
              +xpc10nz) || (6'd52/*MS*/==-8'd64+xpc10nz) || (6'd52/*MS*/==-7'd59+xpc10nz) || (6'd52/*MS*/==-7'd50+xpc10nz) || (6'd52/*MS*/==
              -7'd37+xpc10nz) || (6'd52/*MS*/==-6'd20+xpc10nz) || (6'd52/*MS*/==-6'd19+xpc10nz) || (6'd52/*MS*/==-6'd18+xpc10nz) || (6'd52
              /*MS*/==-6'd17+xpc10nz) || (6'd52/*MS*/==-6'd16+xpc10nz) || (6'd52/*MS*/==-5'd15+xpc10nz) || (6'd52/*MS*/==-5'd14+xpc10nz
              ) || (6'd52/*MS*/==-5'd13+xpc10nz) || (6'd52/*MS*/==-5'd12+xpc10nz) || (6'd52/*MS*/==-5'd11+xpc10nz) || (6'd52/*MS*/==-5'd10
              +xpc10nz) || (6'd52/*MS*/==-5'd9+xpc10nz) || (6'd52/*MS*/==-5'd8+xpc10nz) || (6'd52/*MS*/==-4'd7+xpc10nz) || (6'd52/*MS*/==
              -4'd6+xpc10nz) || (6'd52/*MS*/==-4'd5+xpc10nz) || (6'd52/*MS*/==-4'd4+xpc10nz) || (6'd52/*MS*/==-3'd3+xpc10nz) || (6'd52
              /*MS*/==-3'd2+xpc10nz) || (6'd52/*MS*/==-2'd1+xpc10nz) || (xpc10nz==6'd52/*US*/)) && !xpc10_clear && !xpc10_stall;

               xpc10_trk51 <= ((6'd51/*MS*/==-11'd609+xpc10nz) || (6'd51/*MS*/==-11'd599+xpc10nz) || (6'd51/*MS*/==-11'd588+xpc10nz) || 
              (6'd51/*MS*/==-11'd576+xpc10nz) || (6'd51/*MS*/==-11'd571+xpc10nz) || (6'd51/*MS*/==-11'd565+xpc10nz) || (6'd51/*MS*/==
              -11'd558+xpc10nz) || (6'd51/*MS*/==-11'd550+xpc10nz) || (6'd51/*MS*/==-11'd549+xpc10nz) || (6'd51/*MS*/==-11'd547+xpc10nz
              ) || (6'd51/*MS*/==-11'd544+xpc10nz) || (6'd51/*MS*/==-11'd540+xpc10nz) || (6'd51/*MS*/==-11'd539+xpc10nz) || (6'd51/*MS*/==
              -11'd537+xpc10nz) || (6'd51/*MS*/==-11'd534+xpc10nz) || (6'd51/*MS*/==-11'd532+xpc10nz) || (6'd51/*MS*/==-11'd528+xpc10nz
              ) || (6'd51/*MS*/==-10'd503+xpc10nz) || (6'd51/*MS*/==-10'd502+xpc10nz) || (6'd51/*MS*/==-10'd472+xpc10nz) || (6'd51/*MS*/==
              -10'd407+xpc10nz) || (6'd51/*MS*/==-10'd342+xpc10nz) || (6'd51/*MS*/==-10'd341+xpc10nz) || (6'd51/*MS*/==-10'd340+xpc10nz
              ) || (6'd51/*MS*/==-10'd338+xpc10nz) || (6'd51/*MS*/==-10'd335+xpc10nz) || (6'd51/*MS*/==-10'd334+xpc10nz) || (6'd51/*MS*/==
              -10'd330+xpc10nz) || (6'd51/*MS*/==-10'd329+xpc10nz) || (6'd51/*MS*/==-10'd327+xpc10nz) || (6'd51/*MS*/==-10'd324+xpc10nz
              ) || (6'd51/*MS*/==-10'd323+xpc10nz) || (6'd51/*MS*/==-10'd322+xpc10nz) || (6'd51/*MS*/==-10'd321+xpc10nz) || (6'd51/*MS*/==
              -10'd320+xpc10nz) || (6'd51/*MS*/==-10'd319+xpc10nz) || (6'd51/*MS*/==-10'd318+xpc10nz) || (6'd51/*MS*/==-10'd314+xpc10nz
              ) || (6'd51/*MS*/==-10'd289+xpc10nz) || (6'd51/*MS*/==-10'd287+xpc10nz) || (6'd51/*MS*/==-10'd285+xpc10nz) || (6'd51/*MS*/==
              -10'd284+xpc10nz) || (6'd51/*MS*/==-10'd259+xpc10nz) || (6'd51/*MS*/==-10'd258+xpc10nz) || (6'd51/*MS*/==-10'd257+xpc10nz
              ) || (6'd51/*MS*/==-9'd255+xpc10nz) || (6'd51/*MS*/==-9'd254+xpc10nz) || (6'd51/*MS*/==-9'd253+xpc10nz) || (6'd51/*MS*/==
              -9'd252+xpc10nz) || (6'd51/*MS*/==-9'd251+xpc10nz) || (6'd51/*MS*/==-9'd250+xpc10nz) || (6'd51/*MS*/==-9'd249+xpc10nz) || 
              (6'd51/*MS*/==-9'd248+xpc10nz) || (6'd51/*MS*/==-9'd247+xpc10nz) || (6'd51/*MS*/==-9'd246+xpc10nz) || (6'd51/*MS*/==-9'd245
              +xpc10nz) || (6'd51/*MS*/==-9'd244+xpc10nz) || (6'd51/*MS*/==-9'd242+xpc10nz) || (6'd51/*MS*/==-9'd241+xpc10nz) || (6'd51
              /*MS*/==-9'd239+xpc10nz) || (6'd51/*MS*/==-9'd238+xpc10nz) || (6'd51/*MS*/==-9'd236+xpc10nz) || (6'd51/*MS*/==-9'd171+xpc10nz
              ) || (6'd51/*MS*/==-8'd106+xpc10nz) || (6'd51/*MS*/==-8'd105+xpc10nz) || (6'd51/*MS*/==-8'd104+xpc10nz) || (6'd51/*MS*/==
              -8'd103+xpc10nz) || (6'd51/*MS*/==-8'd102+xpc10nz) || (6'd51/*MS*/==-8'd101+xpc10nz) || (6'd51/*MS*/==-8'd100+xpc10nz) || 
              (6'd51/*MS*/==-8'd99+xpc10nz) || (6'd51/*MS*/==-8'd98+xpc10nz) || (6'd51/*MS*/==-8'd97+xpc10nz) || (6'd51/*MS*/==-8'd96
              +xpc10nz) || (6'd51/*MS*/==-8'd95+xpc10nz) || (6'd51/*MS*/==-8'd94+xpc10nz) || (6'd51/*MS*/==-8'd93+xpc10nz) || (6'd51/*MS*/==
              -8'd92+xpc10nz) || (6'd51/*MS*/==-8'd91+xpc10nz) || (6'd51/*MS*/==-8'd90+xpc10nz) || (6'd51/*MS*/==-8'd89+xpc10nz) || (6'd51
              /*MS*/==-8'd88+xpc10nz) || (6'd51/*MS*/==-8'd87+xpc10nz) || (6'd51/*MS*/==-8'd86+xpc10nz) || (6'd51/*MS*/==-8'd85+xpc10nz
              ) || (6'd51/*MS*/==-8'd84+xpc10nz) || (6'd51/*MS*/==-8'd83+xpc10nz) || (6'd51/*MS*/==-8'd82+xpc10nz) || (6'd51/*MS*/==-8'd65
              +xpc10nz) || (6'd51/*MS*/==-8'd64+xpc10nz) || (6'd51/*MS*/==-7'd59+xpc10nz) || (6'd51/*MS*/==-7'd50+xpc10nz) || (6'd51/*MS*/==
              -7'd37+xpc10nz) || (6'd51/*MS*/==-6'd20+xpc10nz) || (6'd51/*MS*/==-6'd19+xpc10nz) || (6'd51/*MS*/==-6'd18+xpc10nz) || (6'd51
              /*MS*/==-6'd17+xpc10nz) || (6'd51/*MS*/==-6'd16+xpc10nz) || (6'd51/*MS*/==-5'd15+xpc10nz) || (6'd51/*MS*/==-5'd14+xpc10nz
              ) || (6'd51/*MS*/==-5'd13+xpc10nz) || (6'd51/*MS*/==-5'd12+xpc10nz) || (6'd51/*MS*/==-5'd11+xpc10nz) || (6'd51/*MS*/==-5'd10
              +xpc10nz) || (6'd51/*MS*/==-5'd9+xpc10nz) || (6'd51/*MS*/==-5'd8+xpc10nz) || (6'd51/*MS*/==-4'd7+xpc10nz) || (6'd51/*MS*/==
              -4'd6+xpc10nz) || (6'd51/*MS*/==-4'd5+xpc10nz) || (6'd51/*MS*/==-4'd4+xpc10nz) || (6'd51/*MS*/==-3'd3+xpc10nz) || (6'd51
              /*MS*/==-3'd2+xpc10nz) || (6'd51/*MS*/==-2'd1+xpc10nz) || (xpc10nz==6'd51/*US*/)) && !xpc10_clear && !xpc10_stall;

               xpc10_trk50 <= ((6'd50/*MS*/==-11'd609+xpc10nz) || (6'd50/*MS*/==-11'd599+xpc10nz) || (6'd50/*MS*/==-11'd588+xpc10nz) || 
              (6'd50/*MS*/==-11'd576+xpc10nz) || (6'd50/*MS*/==-11'd571+xpc10nz) || (6'd50/*MS*/==-11'd565+xpc10nz) || (6'd50/*MS*/==
              -11'd558+xpc10nz) || (6'd50/*MS*/==-11'd550+xpc10nz) || (6'd50/*MS*/==-11'd549+xpc10nz) || (6'd50/*MS*/==-11'd547+xpc10nz
              ) || (6'd50/*MS*/==-11'd544+xpc10nz) || (6'd50/*MS*/==-11'd540+xpc10nz) || (6'd50/*MS*/==-11'd539+xpc10nz) || (6'd50/*MS*/==
              -11'd537+xpc10nz) || (6'd50/*MS*/==-11'd534+xpc10nz) || (6'd50/*MS*/==-11'd532+xpc10nz) || (6'd50/*MS*/==-11'd528+xpc10nz
              ) || (6'd50/*MS*/==-10'd503+xpc10nz) || (6'd50/*MS*/==-10'd502+xpc10nz) || (6'd50/*MS*/==-10'd472+xpc10nz) || (6'd50/*MS*/==
              -10'd407+xpc10nz) || (6'd50/*MS*/==-10'd342+xpc10nz) || (6'd50/*MS*/==-10'd341+xpc10nz) || (6'd50/*MS*/==-10'd340+xpc10nz
              ) || (6'd50/*MS*/==-10'd338+xpc10nz) || (6'd50/*MS*/==-10'd335+xpc10nz) || (6'd50/*MS*/==-10'd334+xpc10nz) || (6'd50/*MS*/==
              -10'd330+xpc10nz) || (6'd50/*MS*/==-10'd329+xpc10nz) || (6'd50/*MS*/==-10'd327+xpc10nz) || (6'd50/*MS*/==-10'd324+xpc10nz
              ) || (6'd50/*MS*/==-10'd323+xpc10nz) || (6'd50/*MS*/==-10'd322+xpc10nz) || (6'd50/*MS*/==-10'd321+xpc10nz) || (6'd50/*MS*/==
              -10'd320+xpc10nz) || (6'd50/*MS*/==-10'd319+xpc10nz) || (6'd50/*MS*/==-10'd318+xpc10nz) || (6'd50/*MS*/==-10'd314+xpc10nz
              ) || (6'd50/*MS*/==-10'd289+xpc10nz) || (6'd50/*MS*/==-10'd287+xpc10nz) || (6'd50/*MS*/==-10'd285+xpc10nz) || (6'd50/*MS*/==
              -10'd284+xpc10nz) || (6'd50/*MS*/==-10'd259+xpc10nz) || (6'd50/*MS*/==-10'd258+xpc10nz) || (6'd50/*MS*/==-10'd257+xpc10nz
              ) || (6'd50/*MS*/==-9'd255+xpc10nz) || (6'd50/*MS*/==-9'd254+xpc10nz) || (6'd50/*MS*/==-9'd253+xpc10nz) || (6'd50/*MS*/==
              -9'd252+xpc10nz) || (6'd50/*MS*/==-9'd251+xpc10nz) || (6'd50/*MS*/==-9'd250+xpc10nz) || (6'd50/*MS*/==-9'd249+xpc10nz) || 
              (6'd50/*MS*/==-9'd248+xpc10nz) || (6'd50/*MS*/==-9'd247+xpc10nz) || (6'd50/*MS*/==-9'd246+xpc10nz) || (6'd50/*MS*/==-9'd245
              +xpc10nz) || (6'd50/*MS*/==-9'd244+xpc10nz) || (6'd50/*MS*/==-9'd242+xpc10nz) || (6'd50/*MS*/==-9'd241+xpc10nz) || (6'd50
              /*MS*/==-9'd239+xpc10nz) || (6'd50/*MS*/==-9'd238+xpc10nz) || (6'd50/*MS*/==-9'd236+xpc10nz) || (6'd50/*MS*/==-9'd171+xpc10nz
              ) || (6'd50/*MS*/==-8'd106+xpc10nz) || (6'd50/*MS*/==-8'd105+xpc10nz) || (6'd50/*MS*/==-8'd104+xpc10nz) || (6'd50/*MS*/==
              -8'd103+xpc10nz) || (6'd50/*MS*/==-8'd102+xpc10nz) || (6'd50/*MS*/==-8'd101+xpc10nz) || (6'd50/*MS*/==-8'd100+xpc10nz) || 
              (6'd50/*MS*/==-8'd99+xpc10nz) || (6'd50/*MS*/==-8'd98+xpc10nz) || (6'd50/*MS*/==-8'd97+xpc10nz) || (6'd50/*MS*/==-8'd96
              +xpc10nz) || (6'd50/*MS*/==-8'd95+xpc10nz) || (6'd50/*MS*/==-8'd94+xpc10nz) || (6'd50/*MS*/==-8'd93+xpc10nz) || (6'd50/*MS*/==
              -8'd92+xpc10nz) || (6'd50/*MS*/==-8'd91+xpc10nz) || (6'd50/*MS*/==-8'd90+xpc10nz) || (6'd50/*MS*/==-8'd89+xpc10nz) || (6'd50
              /*MS*/==-8'd88+xpc10nz) || (6'd50/*MS*/==-8'd87+xpc10nz) || (6'd50/*MS*/==-8'd86+xpc10nz) || (6'd50/*MS*/==-8'd85+xpc10nz
              ) || (6'd50/*MS*/==-8'd84+xpc10nz) || (6'd50/*MS*/==-8'd83+xpc10nz) || (6'd50/*MS*/==-8'd82+xpc10nz) || (6'd50/*MS*/==-8'd65
              +xpc10nz) || (6'd50/*MS*/==-8'd64+xpc10nz) || (6'd50/*MS*/==-7'd59+xpc10nz) || (6'd50/*MS*/==-7'd50+xpc10nz) || (6'd50/*MS*/==
              -7'd37+xpc10nz) || (6'd50/*MS*/==-6'd20+xpc10nz) || (6'd50/*MS*/==-6'd19+xpc10nz) || (6'd50/*MS*/==-6'd18+xpc10nz) || (6'd50
              /*MS*/==-6'd17+xpc10nz) || (6'd50/*MS*/==-6'd16+xpc10nz) || (6'd50/*MS*/==-5'd15+xpc10nz) || (6'd50/*MS*/==-5'd14+xpc10nz
              ) || (6'd50/*MS*/==-5'd13+xpc10nz) || (6'd50/*MS*/==-5'd12+xpc10nz) || (6'd50/*MS*/==-5'd11+xpc10nz) || (6'd50/*MS*/==-5'd10
              +xpc10nz) || (6'd50/*MS*/==-5'd9+xpc10nz) || (6'd50/*MS*/==-5'd8+xpc10nz) || (6'd50/*MS*/==-4'd7+xpc10nz) || (6'd50/*MS*/==
              -4'd6+xpc10nz) || (6'd50/*MS*/==-4'd5+xpc10nz) || (6'd50/*MS*/==-4'd4+xpc10nz) || (6'd50/*MS*/==-3'd3+xpc10nz) || (6'd50
              /*MS*/==-3'd2+xpc10nz) || (6'd50/*MS*/==-2'd1+xpc10nz) || (xpc10nz==6'd50/*US*/)) && !xpc10_clear && !xpc10_stall;

               xpc10_trk49 <= ((6'd49/*MS*/==-11'd609+xpc10nz) || (6'd49/*MS*/==-11'd599+xpc10nz) || (6'd49/*MS*/==-11'd588+xpc10nz) || 
              (6'd49/*MS*/==-11'd576+xpc10nz) || (6'd49/*MS*/==-11'd571+xpc10nz) || (6'd49/*MS*/==-11'd565+xpc10nz) || (6'd49/*MS*/==
              -11'd558+xpc10nz) || (6'd49/*MS*/==-11'd550+xpc10nz) || (6'd49/*MS*/==-11'd549+xpc10nz) || (6'd49/*MS*/==-11'd547+xpc10nz
              ) || (6'd49/*MS*/==-11'd544+xpc10nz) || (6'd49/*MS*/==-11'd540+xpc10nz) || (6'd49/*MS*/==-11'd539+xpc10nz) || (6'd49/*MS*/==
              -11'd537+xpc10nz) || (6'd49/*MS*/==-11'd534+xpc10nz) || (6'd49/*MS*/==-11'd532+xpc10nz) || (6'd49/*MS*/==-11'd528+xpc10nz
              ) || (6'd49/*MS*/==-10'd503+xpc10nz) || (6'd49/*MS*/==-10'd502+xpc10nz) || (6'd49/*MS*/==-10'd472+xpc10nz) || (6'd49/*MS*/==
              -10'd407+xpc10nz) || (6'd49/*MS*/==-10'd342+xpc10nz) || (6'd49/*MS*/==-10'd341+xpc10nz) || (6'd49/*MS*/==-10'd340+xpc10nz
              ) || (6'd49/*MS*/==-10'd338+xpc10nz) || (6'd49/*MS*/==-10'd335+xpc10nz) || (6'd49/*MS*/==-10'd334+xpc10nz) || (6'd49/*MS*/==
              -10'd330+xpc10nz) || (6'd49/*MS*/==-10'd329+xpc10nz) || (6'd49/*MS*/==-10'd327+xpc10nz) || (6'd49/*MS*/==-10'd324+xpc10nz
              ) || (6'd49/*MS*/==-10'd323+xpc10nz) || (6'd49/*MS*/==-10'd322+xpc10nz) || (6'd49/*MS*/==-10'd321+xpc10nz) || (6'd49/*MS*/==
              -10'd320+xpc10nz) || (6'd49/*MS*/==-10'd319+xpc10nz) || (6'd49/*MS*/==-10'd318+xpc10nz) || (6'd49/*MS*/==-10'd314+xpc10nz
              ) || (6'd49/*MS*/==-10'd289+xpc10nz) || (6'd49/*MS*/==-10'd287+xpc10nz) || (6'd49/*MS*/==-10'd285+xpc10nz) || (6'd49/*MS*/==
              -10'd284+xpc10nz) || (6'd49/*MS*/==-10'd259+xpc10nz) || (6'd49/*MS*/==-10'd258+xpc10nz) || (6'd49/*MS*/==-10'd257+xpc10nz
              ) || (6'd49/*MS*/==-9'd255+xpc10nz) || (6'd49/*MS*/==-9'd254+xpc10nz) || (6'd49/*MS*/==-9'd253+xpc10nz) || (6'd49/*MS*/==
              -9'd252+xpc10nz) || (6'd49/*MS*/==-9'd251+xpc10nz) || (6'd49/*MS*/==-9'd250+xpc10nz) || (6'd49/*MS*/==-9'd249+xpc10nz) || 
              (6'd49/*MS*/==-9'd248+xpc10nz) || (6'd49/*MS*/==-9'd247+xpc10nz) || (6'd49/*MS*/==-9'd246+xpc10nz) || (6'd49/*MS*/==-9'd245
              +xpc10nz) || (6'd49/*MS*/==-9'd244+xpc10nz) || (6'd49/*MS*/==-9'd242+xpc10nz) || (6'd49/*MS*/==-9'd241+xpc10nz) || (6'd49
              /*MS*/==-9'd239+xpc10nz) || (6'd49/*MS*/==-9'd238+xpc10nz) || (6'd49/*MS*/==-9'd236+xpc10nz) || (6'd49/*MS*/==-9'd171+xpc10nz
              ) || (6'd49/*MS*/==-8'd106+xpc10nz) || (6'd49/*MS*/==-8'd105+xpc10nz) || (6'd49/*MS*/==-8'd104+xpc10nz) || (6'd49/*MS*/==
              -8'd103+xpc10nz) || (6'd49/*MS*/==-8'd102+xpc10nz) || (6'd49/*MS*/==-8'd101+xpc10nz) || (6'd49/*MS*/==-8'd100+xpc10nz) || 
              (6'd49/*MS*/==-8'd99+xpc10nz) || (6'd49/*MS*/==-8'd98+xpc10nz) || (6'd49/*MS*/==-8'd97+xpc10nz) || (6'd49/*MS*/==-8'd96
              +xpc10nz) || (6'd49/*MS*/==-8'd95+xpc10nz) || (6'd49/*MS*/==-8'd94+xpc10nz) || (6'd49/*MS*/==-8'd93+xpc10nz) || (6'd49/*MS*/==
              -8'd92+xpc10nz) || (6'd49/*MS*/==-8'd91+xpc10nz) || (6'd49/*MS*/==-8'd90+xpc10nz) || (6'd49/*MS*/==-8'd89+xpc10nz) || (6'd49
              /*MS*/==-8'd88+xpc10nz) || (6'd49/*MS*/==-8'd87+xpc10nz) || (6'd49/*MS*/==-8'd86+xpc10nz) || (6'd49/*MS*/==-8'd85+xpc10nz
              ) || (6'd49/*MS*/==-8'd84+xpc10nz) || (6'd49/*MS*/==-8'd83+xpc10nz) || (6'd49/*MS*/==-8'd82+xpc10nz) || (6'd49/*MS*/==-8'd65
              +xpc10nz) || (6'd49/*MS*/==-8'd64+xpc10nz) || (6'd49/*MS*/==-7'd59+xpc10nz) || (6'd49/*MS*/==-7'd50+xpc10nz) || (6'd49/*MS*/==
              -7'd37+xpc10nz) || (6'd49/*MS*/==-6'd20+xpc10nz) || (6'd49/*MS*/==-6'd19+xpc10nz) || (6'd49/*MS*/==-6'd18+xpc10nz) || (6'd49
              /*MS*/==-6'd17+xpc10nz) || (6'd49/*MS*/==-6'd16+xpc10nz) || (6'd49/*MS*/==-5'd15+xpc10nz) || (6'd49/*MS*/==-5'd14+xpc10nz
              ) || (6'd49/*MS*/==-5'd13+xpc10nz) || (6'd49/*MS*/==-5'd12+xpc10nz) || (6'd49/*MS*/==-5'd11+xpc10nz) || (6'd49/*MS*/==-5'd10
              +xpc10nz) || (6'd49/*MS*/==-5'd9+xpc10nz) || (6'd49/*MS*/==-5'd8+xpc10nz) || (6'd49/*MS*/==-4'd7+xpc10nz) || (6'd49/*MS*/==
              -4'd6+xpc10nz) || (6'd49/*MS*/==-4'd5+xpc10nz) || (6'd49/*MS*/==-4'd4+xpc10nz) || (6'd49/*MS*/==-3'd3+xpc10nz) || (6'd49
              /*MS*/==-3'd2+xpc10nz) || (6'd49/*MS*/==-2'd1+xpc10nz) || (xpc10nz==6'd49/*US*/)) && !xpc10_clear && !xpc10_stall;

               xpc10_trk48 <= ((6'd48/*MS*/==-11'd609+xpc10nz) || (6'd48/*MS*/==-11'd599+xpc10nz) || (6'd48/*MS*/==-11'd588+xpc10nz) || 
              (6'd48/*MS*/==-11'd576+xpc10nz) || (6'd48/*MS*/==-11'd571+xpc10nz) || (6'd48/*MS*/==-11'd565+xpc10nz) || (6'd48/*MS*/==
              -11'd558+xpc10nz) || (6'd48/*MS*/==-11'd550+xpc10nz) || (6'd48/*MS*/==-11'd549+xpc10nz) || (6'd48/*MS*/==-11'd547+xpc10nz
              ) || (6'd48/*MS*/==-11'd544+xpc10nz) || (6'd48/*MS*/==-11'd540+xpc10nz) || (6'd48/*MS*/==-11'd539+xpc10nz) || (6'd48/*MS*/==
              -11'd537+xpc10nz) || (6'd48/*MS*/==-11'd534+xpc10nz) || (6'd48/*MS*/==-11'd532+xpc10nz) || (6'd48/*MS*/==-11'd528+xpc10nz
              ) || (6'd48/*MS*/==-10'd503+xpc10nz) || (6'd48/*MS*/==-10'd502+xpc10nz) || (6'd48/*MS*/==-10'd472+xpc10nz) || (6'd48/*MS*/==
              -10'd407+xpc10nz) || (6'd48/*MS*/==-10'd342+xpc10nz) || (6'd48/*MS*/==-10'd341+xpc10nz) || (6'd48/*MS*/==-10'd340+xpc10nz
              ) || (6'd48/*MS*/==-10'd338+xpc10nz) || (6'd48/*MS*/==-10'd335+xpc10nz) || (6'd48/*MS*/==-10'd334+xpc10nz) || (6'd48/*MS*/==
              -10'd330+xpc10nz) || (6'd48/*MS*/==-10'd329+xpc10nz) || (6'd48/*MS*/==-10'd327+xpc10nz) || (6'd48/*MS*/==-10'd324+xpc10nz
              ) || (6'd48/*MS*/==-10'd323+xpc10nz) || (6'd48/*MS*/==-10'd322+xpc10nz) || (6'd48/*MS*/==-10'd321+xpc10nz) || (6'd48/*MS*/==
              -10'd320+xpc10nz) || (6'd48/*MS*/==-10'd319+xpc10nz) || (6'd48/*MS*/==-10'd318+xpc10nz) || (6'd48/*MS*/==-10'd314+xpc10nz
              ) || (6'd48/*MS*/==-10'd289+xpc10nz) || (6'd48/*MS*/==-10'd287+xpc10nz) || (6'd48/*MS*/==-10'd285+xpc10nz) || (6'd48/*MS*/==
              -10'd284+xpc10nz) || (6'd48/*MS*/==-10'd259+xpc10nz) || (6'd48/*MS*/==-10'd258+xpc10nz) || (6'd48/*MS*/==-10'd257+xpc10nz
              ) || (6'd48/*MS*/==-9'd255+xpc10nz) || (6'd48/*MS*/==-9'd254+xpc10nz) || (6'd48/*MS*/==-9'd253+xpc10nz) || (6'd48/*MS*/==
              -9'd252+xpc10nz) || (6'd48/*MS*/==-9'd251+xpc10nz) || (6'd48/*MS*/==-9'd250+xpc10nz) || (6'd48/*MS*/==-9'd249+xpc10nz) || 
              (6'd48/*MS*/==-9'd248+xpc10nz) || (6'd48/*MS*/==-9'd247+xpc10nz) || (6'd48/*MS*/==-9'd246+xpc10nz) || (6'd48/*MS*/==-9'd245
              +xpc10nz) || (6'd48/*MS*/==-9'd244+xpc10nz) || (6'd48/*MS*/==-9'd242+xpc10nz) || (6'd48/*MS*/==-9'd241+xpc10nz) || (6'd48
              /*MS*/==-9'd239+xpc10nz) || (6'd48/*MS*/==-9'd238+xpc10nz) || (6'd48/*MS*/==-9'd236+xpc10nz) || (6'd48/*MS*/==-9'd171+xpc10nz
              ) || (6'd48/*MS*/==-8'd106+xpc10nz) || (6'd48/*MS*/==-8'd105+xpc10nz) || (6'd48/*MS*/==-8'd104+xpc10nz) || (6'd48/*MS*/==
              -8'd103+xpc10nz) || (6'd48/*MS*/==-8'd102+xpc10nz) || (6'd48/*MS*/==-8'd101+xpc10nz) || (6'd48/*MS*/==-8'd100+xpc10nz) || 
              (6'd48/*MS*/==-8'd99+xpc10nz) || (6'd48/*MS*/==-8'd98+xpc10nz) || (6'd48/*MS*/==-8'd97+xpc10nz) || (6'd48/*MS*/==-8'd96
              +xpc10nz) || (6'd48/*MS*/==-8'd95+xpc10nz) || (6'd48/*MS*/==-8'd94+xpc10nz) || (6'd48/*MS*/==-8'd93+xpc10nz) || (6'd48/*MS*/==
              -8'd92+xpc10nz) || (6'd48/*MS*/==-8'd91+xpc10nz) || (6'd48/*MS*/==-8'd90+xpc10nz) || (6'd48/*MS*/==-8'd89+xpc10nz) || (6'd48
              /*MS*/==-8'd88+xpc10nz) || (6'd48/*MS*/==-8'd87+xpc10nz) || (6'd48/*MS*/==-8'd86+xpc10nz) || (6'd48/*MS*/==-8'd85+xpc10nz
              ) || (6'd48/*MS*/==-8'd84+xpc10nz) || (6'd48/*MS*/==-8'd83+xpc10nz) || (6'd48/*MS*/==-8'd82+xpc10nz) || (6'd48/*MS*/==-8'd65
              +xpc10nz) || (6'd48/*MS*/==-8'd64+xpc10nz) || (6'd48/*MS*/==-7'd59+xpc10nz) || (6'd48/*MS*/==-7'd50+xpc10nz) || (6'd48/*MS*/==
              -7'd37+xpc10nz) || (6'd48/*MS*/==-6'd20+xpc10nz) || (6'd48/*MS*/==-6'd19+xpc10nz) || (6'd48/*MS*/==-6'd18+xpc10nz) || (6'd48
              /*MS*/==-6'd17+xpc10nz) || (6'd48/*MS*/==-6'd16+xpc10nz) || (6'd48/*MS*/==-5'd15+xpc10nz) || (6'd48/*MS*/==-5'd14+xpc10nz
              ) || (6'd48/*MS*/==-5'd13+xpc10nz) || (6'd48/*MS*/==-5'd12+xpc10nz) || (6'd48/*MS*/==-5'd11+xpc10nz) || (6'd48/*MS*/==-5'd10
              +xpc10nz) || (6'd48/*MS*/==-5'd9+xpc10nz) || (6'd48/*MS*/==-5'd8+xpc10nz) || (6'd48/*MS*/==-4'd7+xpc10nz) || (6'd48/*MS*/==
              -4'd6+xpc10nz) || (6'd48/*MS*/==-4'd5+xpc10nz) || (6'd48/*MS*/==-4'd4+xpc10nz) || (6'd48/*MS*/==-3'd3+xpc10nz) || (6'd48
              /*MS*/==-3'd2+xpc10nz) || (6'd48/*MS*/==-2'd1+xpc10nz) || (xpc10nz==6'd48/*US*/)) && !xpc10_clear && !xpc10_stall;

               xpc10_trk47 <= ((6'd47/*MS*/==-11'd609+xpc10nz) || (6'd47/*MS*/==-11'd599+xpc10nz) || (6'd47/*MS*/==-11'd588+xpc10nz) || 
              (6'd47/*MS*/==-11'd576+xpc10nz) || (6'd47/*MS*/==-11'd571+xpc10nz) || (6'd47/*MS*/==-11'd565+xpc10nz) || (6'd47/*MS*/==
              -11'd558+xpc10nz) || (6'd47/*MS*/==-11'd550+xpc10nz) || (6'd47/*MS*/==-11'd549+xpc10nz) || (6'd47/*MS*/==-11'd547+xpc10nz
              ) || (6'd47/*MS*/==-11'd544+xpc10nz) || (6'd47/*MS*/==-11'd540+xpc10nz) || (6'd47/*MS*/==-11'd539+xpc10nz) || (6'd47/*MS*/==
              -11'd537+xpc10nz) || (6'd47/*MS*/==-11'd534+xpc10nz) || (6'd47/*MS*/==-11'd532+xpc10nz) || (6'd47/*MS*/==-11'd528+xpc10nz
              ) || (6'd47/*MS*/==-10'd503+xpc10nz) || (6'd47/*MS*/==-10'd502+xpc10nz) || (6'd47/*MS*/==-10'd472+xpc10nz) || (6'd47/*MS*/==
              -10'd407+xpc10nz) || (6'd47/*MS*/==-10'd342+xpc10nz) || (6'd47/*MS*/==-10'd341+xpc10nz) || (6'd47/*MS*/==-10'd340+xpc10nz
              ) || (6'd47/*MS*/==-10'd338+xpc10nz) || (6'd47/*MS*/==-10'd335+xpc10nz) || (6'd47/*MS*/==-10'd334+xpc10nz) || (6'd47/*MS*/==
              -10'd330+xpc10nz) || (6'd47/*MS*/==-10'd329+xpc10nz) || (6'd47/*MS*/==-10'd327+xpc10nz) || (6'd47/*MS*/==-10'd324+xpc10nz
              ) || (6'd47/*MS*/==-10'd323+xpc10nz) || (6'd47/*MS*/==-10'd322+xpc10nz) || (6'd47/*MS*/==-10'd321+xpc10nz) || (6'd47/*MS*/==
              -10'd320+xpc10nz) || (6'd47/*MS*/==-10'd319+xpc10nz) || (6'd47/*MS*/==-10'd318+xpc10nz) || (6'd47/*MS*/==-10'd314+xpc10nz
              ) || (6'd47/*MS*/==-10'd289+xpc10nz) || (6'd47/*MS*/==-10'd287+xpc10nz) || (6'd47/*MS*/==-10'd285+xpc10nz) || (6'd47/*MS*/==
              -10'd284+xpc10nz) || (6'd47/*MS*/==-10'd259+xpc10nz) || (6'd47/*MS*/==-10'd258+xpc10nz) || (6'd47/*MS*/==-10'd257+xpc10nz
              ) || (6'd47/*MS*/==-9'd255+xpc10nz) || (6'd47/*MS*/==-9'd254+xpc10nz) || (6'd47/*MS*/==-9'd253+xpc10nz) || (6'd47/*MS*/==
              -9'd252+xpc10nz) || (6'd47/*MS*/==-9'd251+xpc10nz) || (6'd47/*MS*/==-9'd250+xpc10nz) || (6'd47/*MS*/==-9'd249+xpc10nz) || 
              (6'd47/*MS*/==-9'd248+xpc10nz) || (6'd47/*MS*/==-9'd247+xpc10nz) || (6'd47/*MS*/==-9'd246+xpc10nz) || (6'd47/*MS*/==-9'd245
              +xpc10nz) || (6'd47/*MS*/==-9'd244+xpc10nz) || (6'd47/*MS*/==-9'd242+xpc10nz) || (6'd47/*MS*/==-9'd241+xpc10nz) || (6'd47
              /*MS*/==-9'd239+xpc10nz) || (6'd47/*MS*/==-9'd238+xpc10nz) || (6'd47/*MS*/==-9'd236+xpc10nz) || (6'd47/*MS*/==-9'd171+xpc10nz
              ) || (6'd47/*MS*/==-8'd106+xpc10nz) || (6'd47/*MS*/==-8'd105+xpc10nz) || (6'd47/*MS*/==-8'd104+xpc10nz) || (6'd47/*MS*/==
              -8'd103+xpc10nz) || (6'd47/*MS*/==-8'd102+xpc10nz) || (6'd47/*MS*/==-8'd101+xpc10nz) || (6'd47/*MS*/==-8'd100+xpc10nz) || 
              (6'd47/*MS*/==-8'd99+xpc10nz) || (6'd47/*MS*/==-8'd98+xpc10nz) || (6'd47/*MS*/==-8'd97+xpc10nz) || (6'd47/*MS*/==-8'd96
              +xpc10nz) || (6'd47/*MS*/==-8'd95+xpc10nz) || (6'd47/*MS*/==-8'd94+xpc10nz) || (6'd47/*MS*/==-8'd93+xpc10nz) || (6'd47/*MS*/==
              -8'd92+xpc10nz) || (6'd47/*MS*/==-8'd91+xpc10nz) || (6'd47/*MS*/==-8'd90+xpc10nz) || (6'd47/*MS*/==-8'd89+xpc10nz) || (6'd47
              /*MS*/==-8'd88+xpc10nz) || (6'd47/*MS*/==-8'd87+xpc10nz) || (6'd47/*MS*/==-8'd86+xpc10nz) || (6'd47/*MS*/==-8'd85+xpc10nz
              ) || (6'd47/*MS*/==-8'd84+xpc10nz) || (6'd47/*MS*/==-8'd83+xpc10nz) || (6'd47/*MS*/==-8'd82+xpc10nz) || (6'd47/*MS*/==-8'd65
              +xpc10nz) || (6'd47/*MS*/==-8'd64+xpc10nz) || (6'd47/*MS*/==-7'd59+xpc10nz) || (6'd47/*MS*/==-7'd50+xpc10nz) || (6'd47/*MS*/==
              -7'd37+xpc10nz) || (6'd47/*MS*/==-6'd20+xpc10nz) || (6'd47/*MS*/==-6'd19+xpc10nz) || (6'd47/*MS*/==-6'd18+xpc10nz) || (6'd47
              /*MS*/==-6'd17+xpc10nz) || (6'd47/*MS*/==-6'd16+xpc10nz) || (6'd47/*MS*/==-5'd15+xpc10nz) || (6'd47/*MS*/==-5'd14+xpc10nz
              ) || (6'd47/*MS*/==-5'd13+xpc10nz) || (6'd47/*MS*/==-5'd12+xpc10nz) || (6'd47/*MS*/==-5'd11+xpc10nz) || (6'd47/*MS*/==-5'd10
              +xpc10nz) || (6'd47/*MS*/==-5'd9+xpc10nz) || (6'd47/*MS*/==-5'd8+xpc10nz) || (6'd47/*MS*/==-4'd7+xpc10nz) || (6'd47/*MS*/==
              -4'd6+xpc10nz) || (6'd47/*MS*/==-4'd5+xpc10nz) || (6'd47/*MS*/==-4'd4+xpc10nz) || (6'd47/*MS*/==-3'd3+xpc10nz) || (6'd47
              /*MS*/==-3'd2+xpc10nz) || (6'd47/*MS*/==-2'd1+xpc10nz) || (xpc10nz==6'd47/*US*/)) && !xpc10_clear && !xpc10_stall;

               xpc10_trk46 <= ((6'd46/*MS*/==-11'd609+xpc10nz) || (6'd46/*MS*/==-11'd599+xpc10nz) || (6'd46/*MS*/==-11'd588+xpc10nz) || 
              (6'd46/*MS*/==-11'd576+xpc10nz) || (6'd46/*MS*/==-11'd571+xpc10nz) || (6'd46/*MS*/==-11'd565+xpc10nz) || (6'd46/*MS*/==
              -11'd558+xpc10nz) || (6'd46/*MS*/==-11'd550+xpc10nz) || (6'd46/*MS*/==-11'd549+xpc10nz) || (6'd46/*MS*/==-11'd547+xpc10nz
              ) || (6'd46/*MS*/==-11'd544+xpc10nz) || (6'd46/*MS*/==-11'd540+xpc10nz) || (6'd46/*MS*/==-11'd539+xpc10nz) || (6'd46/*MS*/==
              -11'd537+xpc10nz) || (6'd46/*MS*/==-11'd534+xpc10nz) || (6'd46/*MS*/==-11'd532+xpc10nz) || (6'd46/*MS*/==-11'd528+xpc10nz
              ) || (6'd46/*MS*/==-10'd503+xpc10nz) || (6'd46/*MS*/==-10'd502+xpc10nz) || (6'd46/*MS*/==-10'd472+xpc10nz) || (6'd46/*MS*/==
              -10'd407+xpc10nz) || (6'd46/*MS*/==-10'd342+xpc10nz) || (6'd46/*MS*/==-10'd341+xpc10nz) || (6'd46/*MS*/==-10'd340+xpc10nz
              ) || (6'd46/*MS*/==-10'd338+xpc10nz) || (6'd46/*MS*/==-10'd335+xpc10nz) || (6'd46/*MS*/==-10'd334+xpc10nz) || (6'd46/*MS*/==
              -10'd330+xpc10nz) || (6'd46/*MS*/==-10'd329+xpc10nz) || (6'd46/*MS*/==-10'd327+xpc10nz) || (6'd46/*MS*/==-10'd324+xpc10nz
              ) || (6'd46/*MS*/==-10'd323+xpc10nz) || (6'd46/*MS*/==-10'd322+xpc10nz) || (6'd46/*MS*/==-10'd321+xpc10nz) || (6'd46/*MS*/==
              -10'd320+xpc10nz) || (6'd46/*MS*/==-10'd319+xpc10nz) || (6'd46/*MS*/==-10'd318+xpc10nz) || (6'd46/*MS*/==-10'd314+xpc10nz
              ) || (6'd46/*MS*/==-10'd289+xpc10nz) || (6'd46/*MS*/==-10'd287+xpc10nz) || (6'd46/*MS*/==-10'd285+xpc10nz) || (6'd46/*MS*/==
              -10'd284+xpc10nz) || (6'd46/*MS*/==-10'd259+xpc10nz) || (6'd46/*MS*/==-10'd258+xpc10nz) || (6'd46/*MS*/==-10'd257+xpc10nz
              ) || (6'd46/*MS*/==-9'd255+xpc10nz) || (6'd46/*MS*/==-9'd254+xpc10nz) || (6'd46/*MS*/==-9'd253+xpc10nz) || (6'd46/*MS*/==
              -9'd252+xpc10nz) || (6'd46/*MS*/==-9'd251+xpc10nz) || (6'd46/*MS*/==-9'd250+xpc10nz) || (6'd46/*MS*/==-9'd249+xpc10nz) || 
              (6'd46/*MS*/==-9'd248+xpc10nz) || (6'd46/*MS*/==-9'd247+xpc10nz) || (6'd46/*MS*/==-9'd246+xpc10nz) || (6'd46/*MS*/==-9'd245
              +xpc10nz) || (6'd46/*MS*/==-9'd244+xpc10nz) || (6'd46/*MS*/==-9'd242+xpc10nz) || (6'd46/*MS*/==-9'd241+xpc10nz) || (6'd46
              /*MS*/==-9'd239+xpc10nz) || (6'd46/*MS*/==-9'd238+xpc10nz) || (6'd46/*MS*/==-9'd236+xpc10nz) || (6'd46/*MS*/==-9'd171+xpc10nz
              ) || (6'd46/*MS*/==-8'd106+xpc10nz) || (6'd46/*MS*/==-8'd105+xpc10nz) || (6'd46/*MS*/==-8'd104+xpc10nz) || (6'd46/*MS*/==
              -8'd103+xpc10nz) || (6'd46/*MS*/==-8'd102+xpc10nz) || (6'd46/*MS*/==-8'd101+xpc10nz) || (6'd46/*MS*/==-8'd100+xpc10nz) || 
              (6'd46/*MS*/==-8'd99+xpc10nz) || (6'd46/*MS*/==-8'd98+xpc10nz) || (6'd46/*MS*/==-8'd97+xpc10nz) || (6'd46/*MS*/==-8'd96
              +xpc10nz) || (6'd46/*MS*/==-8'd95+xpc10nz) || (6'd46/*MS*/==-8'd94+xpc10nz) || (6'd46/*MS*/==-8'd93+xpc10nz) || (6'd46/*MS*/==
              -8'd92+xpc10nz) || (6'd46/*MS*/==-8'd91+xpc10nz) || (6'd46/*MS*/==-8'd90+xpc10nz) || (6'd46/*MS*/==-8'd89+xpc10nz) || (6'd46
              /*MS*/==-8'd88+xpc10nz) || (6'd46/*MS*/==-8'd87+xpc10nz) || (6'd46/*MS*/==-8'd86+xpc10nz) || (6'd46/*MS*/==-8'd85+xpc10nz
              ) || (6'd46/*MS*/==-8'd84+xpc10nz) || (6'd46/*MS*/==-8'd83+xpc10nz) || (6'd46/*MS*/==-8'd82+xpc10nz) || (6'd46/*MS*/==-8'd65
              +xpc10nz) || (6'd46/*MS*/==-8'd64+xpc10nz) || (6'd46/*MS*/==-7'd59+xpc10nz) || (6'd46/*MS*/==-7'd50+xpc10nz) || (6'd46/*MS*/==
              -7'd37+xpc10nz) || (6'd46/*MS*/==-6'd20+xpc10nz) || (6'd46/*MS*/==-6'd19+xpc10nz) || (6'd46/*MS*/==-6'd18+xpc10nz) || (6'd46
              /*MS*/==-6'd17+xpc10nz) || (6'd46/*MS*/==-6'd16+xpc10nz) || (6'd46/*MS*/==-5'd15+xpc10nz) || (6'd46/*MS*/==-5'd14+xpc10nz
              ) || (6'd46/*MS*/==-5'd13+xpc10nz) || (6'd46/*MS*/==-5'd12+xpc10nz) || (6'd46/*MS*/==-5'd11+xpc10nz) || (6'd46/*MS*/==-5'd10
              +xpc10nz) || (6'd46/*MS*/==-5'd9+xpc10nz) || (6'd46/*MS*/==-5'd8+xpc10nz) || (6'd46/*MS*/==-4'd7+xpc10nz) || (6'd46/*MS*/==
              -4'd6+xpc10nz) || (6'd46/*MS*/==-4'd5+xpc10nz) || (6'd46/*MS*/==-4'd4+xpc10nz) || (6'd46/*MS*/==-3'd3+xpc10nz) || (6'd46
              /*MS*/==-3'd2+xpc10nz) || (6'd46/*MS*/==-2'd1+xpc10nz) || (xpc10nz==6'd46/*US*/)) && !xpc10_clear && !xpc10_stall;

               xpc10_trk45 <= ((6'd45/*MS*/==-11'd609+xpc10nz) || (6'd45/*MS*/==-11'd599+xpc10nz) || (6'd45/*MS*/==-11'd588+xpc10nz) || 
              (6'd45/*MS*/==-11'd576+xpc10nz) || (6'd45/*MS*/==-11'd571+xpc10nz) || (6'd45/*MS*/==-11'd565+xpc10nz) || (6'd45/*MS*/==
              -11'd558+xpc10nz) || (6'd45/*MS*/==-11'd550+xpc10nz) || (6'd45/*MS*/==-11'd549+xpc10nz) || (6'd45/*MS*/==-11'd547+xpc10nz
              ) || (6'd45/*MS*/==-11'd544+xpc10nz) || (6'd45/*MS*/==-11'd540+xpc10nz) || (6'd45/*MS*/==-11'd539+xpc10nz) || (6'd45/*MS*/==
              -11'd537+xpc10nz) || (6'd45/*MS*/==-11'd534+xpc10nz) || (6'd45/*MS*/==-11'd532+xpc10nz) || (6'd45/*MS*/==-11'd528+xpc10nz
              ) || (6'd45/*MS*/==-10'd503+xpc10nz) || (6'd45/*MS*/==-10'd502+xpc10nz) || (6'd45/*MS*/==-10'd472+xpc10nz) || (6'd45/*MS*/==
              -10'd407+xpc10nz) || (6'd45/*MS*/==-10'd342+xpc10nz) || (6'd45/*MS*/==-10'd341+xpc10nz) || (6'd45/*MS*/==-10'd340+xpc10nz
              ) || (6'd45/*MS*/==-10'd338+xpc10nz) || (6'd45/*MS*/==-10'd335+xpc10nz) || (6'd45/*MS*/==-10'd334+xpc10nz) || (6'd45/*MS*/==
              -10'd330+xpc10nz) || (6'd45/*MS*/==-10'd329+xpc10nz) || (6'd45/*MS*/==-10'd327+xpc10nz) || (6'd45/*MS*/==-10'd324+xpc10nz
              ) || (6'd45/*MS*/==-10'd323+xpc10nz) || (6'd45/*MS*/==-10'd322+xpc10nz) || (6'd45/*MS*/==-10'd321+xpc10nz) || (6'd45/*MS*/==
              -10'd320+xpc10nz) || (6'd45/*MS*/==-10'd319+xpc10nz) || (6'd45/*MS*/==-10'd318+xpc10nz) || (6'd45/*MS*/==-10'd314+xpc10nz
              ) || (6'd45/*MS*/==-10'd289+xpc10nz) || (6'd45/*MS*/==-10'd287+xpc10nz) || (6'd45/*MS*/==-10'd285+xpc10nz) || (6'd45/*MS*/==
              -10'd284+xpc10nz) || (6'd45/*MS*/==-10'd259+xpc10nz) || (6'd45/*MS*/==-10'd258+xpc10nz) || (6'd45/*MS*/==-10'd257+xpc10nz
              ) || (6'd45/*MS*/==-9'd255+xpc10nz) || (6'd45/*MS*/==-9'd254+xpc10nz) || (6'd45/*MS*/==-9'd253+xpc10nz) || (6'd45/*MS*/==
              -9'd252+xpc10nz) || (6'd45/*MS*/==-9'd251+xpc10nz) || (6'd45/*MS*/==-9'd250+xpc10nz) || (6'd45/*MS*/==-9'd249+xpc10nz) || 
              (6'd45/*MS*/==-9'd248+xpc10nz) || (6'd45/*MS*/==-9'd247+xpc10nz) || (6'd45/*MS*/==-9'd246+xpc10nz) || (6'd45/*MS*/==-9'd245
              +xpc10nz) || (6'd45/*MS*/==-9'd244+xpc10nz) || (6'd45/*MS*/==-9'd242+xpc10nz) || (6'd45/*MS*/==-9'd241+xpc10nz) || (6'd45
              /*MS*/==-9'd239+xpc10nz) || (6'd45/*MS*/==-9'd238+xpc10nz) || (6'd45/*MS*/==-9'd236+xpc10nz) || (6'd45/*MS*/==-9'd171+xpc10nz
              ) || (6'd45/*MS*/==-8'd106+xpc10nz) || (6'd45/*MS*/==-8'd105+xpc10nz) || (6'd45/*MS*/==-8'd104+xpc10nz) || (6'd45/*MS*/==
              -8'd103+xpc10nz) || (6'd45/*MS*/==-8'd102+xpc10nz) || (6'd45/*MS*/==-8'd101+xpc10nz) || (6'd45/*MS*/==-8'd100+xpc10nz) || 
              (6'd45/*MS*/==-8'd99+xpc10nz) || (6'd45/*MS*/==-8'd98+xpc10nz) || (6'd45/*MS*/==-8'd97+xpc10nz) || (6'd45/*MS*/==-8'd96
              +xpc10nz) || (6'd45/*MS*/==-8'd95+xpc10nz) || (6'd45/*MS*/==-8'd94+xpc10nz) || (6'd45/*MS*/==-8'd93+xpc10nz) || (6'd45/*MS*/==
              -8'd92+xpc10nz) || (6'd45/*MS*/==-8'd91+xpc10nz) || (6'd45/*MS*/==-8'd90+xpc10nz) || (6'd45/*MS*/==-8'd89+xpc10nz) || (6'd45
              /*MS*/==-8'd88+xpc10nz) || (6'd45/*MS*/==-8'd87+xpc10nz) || (6'd45/*MS*/==-8'd86+xpc10nz) || (6'd45/*MS*/==-8'd85+xpc10nz
              ) || (6'd45/*MS*/==-8'd84+xpc10nz) || (6'd45/*MS*/==-8'd83+xpc10nz) || (6'd45/*MS*/==-8'd82+xpc10nz) || (6'd45/*MS*/==-8'd65
              +xpc10nz) || (6'd45/*MS*/==-8'd64+xpc10nz) || (6'd45/*MS*/==-7'd59+xpc10nz) || (6'd45/*MS*/==-7'd50+xpc10nz) || (6'd45/*MS*/==
              -7'd37+xpc10nz) || (6'd45/*MS*/==-6'd20+xpc10nz) || (6'd45/*MS*/==-6'd19+xpc10nz) || (6'd45/*MS*/==-6'd18+xpc10nz) || (6'd45
              /*MS*/==-6'd17+xpc10nz) || (6'd45/*MS*/==-6'd16+xpc10nz) || (6'd45/*MS*/==-5'd15+xpc10nz) || (6'd45/*MS*/==-5'd14+xpc10nz
              ) || (6'd45/*MS*/==-5'd13+xpc10nz) || (6'd45/*MS*/==-5'd12+xpc10nz) || (6'd45/*MS*/==-5'd11+xpc10nz) || (6'd45/*MS*/==-5'd10
              +xpc10nz) || (6'd45/*MS*/==-5'd9+xpc10nz) || (6'd45/*MS*/==-5'd8+xpc10nz) || (6'd45/*MS*/==-4'd7+xpc10nz) || (6'd45/*MS*/==
              -4'd6+xpc10nz) || (6'd45/*MS*/==-4'd5+xpc10nz) || (6'd45/*MS*/==-4'd4+xpc10nz) || (6'd45/*MS*/==-3'd3+xpc10nz) || (6'd45
              /*MS*/==-3'd2+xpc10nz) || (6'd45/*MS*/==-2'd1+xpc10nz) || (xpc10nz==6'd45/*US*/)) && !xpc10_clear && !xpc10_stall;

               xpc10_trk44 <= ((6'd44/*MS*/==-11'd609+xpc10nz) || (6'd44/*MS*/==-11'd599+xpc10nz) || (6'd44/*MS*/==-11'd588+xpc10nz) || 
              (6'd44/*MS*/==-11'd576+xpc10nz) || (6'd44/*MS*/==-11'd571+xpc10nz) || (6'd44/*MS*/==-11'd565+xpc10nz) || (6'd44/*MS*/==
              -11'd558+xpc10nz) || (6'd44/*MS*/==-11'd550+xpc10nz) || (6'd44/*MS*/==-11'd549+xpc10nz) || (6'd44/*MS*/==-11'd547+xpc10nz
              ) || (6'd44/*MS*/==-11'd544+xpc10nz) || (6'd44/*MS*/==-11'd540+xpc10nz) || (6'd44/*MS*/==-11'd539+xpc10nz) || (6'd44/*MS*/==
              -11'd537+xpc10nz) || (6'd44/*MS*/==-11'd534+xpc10nz) || (6'd44/*MS*/==-11'd532+xpc10nz) || (6'd44/*MS*/==-11'd528+xpc10nz
              ) || (6'd44/*MS*/==-10'd503+xpc10nz) || (6'd44/*MS*/==-10'd502+xpc10nz) || (6'd44/*MS*/==-10'd472+xpc10nz) || (6'd44/*MS*/==
              -10'd407+xpc10nz) || (6'd44/*MS*/==-10'd342+xpc10nz) || (6'd44/*MS*/==-10'd341+xpc10nz) || (6'd44/*MS*/==-10'd340+xpc10nz
              ) || (6'd44/*MS*/==-10'd338+xpc10nz) || (6'd44/*MS*/==-10'd335+xpc10nz) || (6'd44/*MS*/==-10'd334+xpc10nz) || (6'd44/*MS*/==
              -10'd330+xpc10nz) || (6'd44/*MS*/==-10'd329+xpc10nz) || (6'd44/*MS*/==-10'd327+xpc10nz) || (6'd44/*MS*/==-10'd324+xpc10nz
              ) || (6'd44/*MS*/==-10'd323+xpc10nz) || (6'd44/*MS*/==-10'd322+xpc10nz) || (6'd44/*MS*/==-10'd321+xpc10nz) || (6'd44/*MS*/==
              -10'd320+xpc10nz) || (6'd44/*MS*/==-10'd319+xpc10nz) || (6'd44/*MS*/==-10'd318+xpc10nz) || (6'd44/*MS*/==-10'd314+xpc10nz
              ) || (6'd44/*MS*/==-10'd289+xpc10nz) || (6'd44/*MS*/==-10'd287+xpc10nz) || (6'd44/*MS*/==-10'd285+xpc10nz) || (6'd44/*MS*/==
              -10'd284+xpc10nz) || (6'd44/*MS*/==-10'd259+xpc10nz) || (6'd44/*MS*/==-10'd258+xpc10nz) || (6'd44/*MS*/==-10'd257+xpc10nz
              ) || (6'd44/*MS*/==-9'd255+xpc10nz) || (6'd44/*MS*/==-9'd254+xpc10nz) || (6'd44/*MS*/==-9'd253+xpc10nz) || (6'd44/*MS*/==
              -9'd252+xpc10nz) || (6'd44/*MS*/==-9'd251+xpc10nz) || (6'd44/*MS*/==-9'd250+xpc10nz) || (6'd44/*MS*/==-9'd249+xpc10nz) || 
              (6'd44/*MS*/==-9'd248+xpc10nz) || (6'd44/*MS*/==-9'd247+xpc10nz) || (6'd44/*MS*/==-9'd246+xpc10nz) || (6'd44/*MS*/==-9'd245
              +xpc10nz) || (6'd44/*MS*/==-9'd244+xpc10nz) || (6'd44/*MS*/==-9'd242+xpc10nz) || (6'd44/*MS*/==-9'd241+xpc10nz) || (6'd44
              /*MS*/==-9'd239+xpc10nz) || (6'd44/*MS*/==-9'd238+xpc10nz) || (6'd44/*MS*/==-9'd236+xpc10nz) || (6'd44/*MS*/==-9'd171+xpc10nz
              ) || (6'd44/*MS*/==-8'd106+xpc10nz) || (6'd44/*MS*/==-8'd105+xpc10nz) || (6'd44/*MS*/==-8'd104+xpc10nz) || (6'd44/*MS*/==
              -8'd103+xpc10nz) || (6'd44/*MS*/==-8'd102+xpc10nz) || (6'd44/*MS*/==-8'd101+xpc10nz) || (6'd44/*MS*/==-8'd100+xpc10nz) || 
              (6'd44/*MS*/==-8'd99+xpc10nz) || (6'd44/*MS*/==-8'd98+xpc10nz) || (6'd44/*MS*/==-8'd97+xpc10nz) || (6'd44/*MS*/==-8'd96
              +xpc10nz) || (6'd44/*MS*/==-8'd95+xpc10nz) || (6'd44/*MS*/==-8'd94+xpc10nz) || (6'd44/*MS*/==-8'd93+xpc10nz) || (6'd44/*MS*/==
              -8'd92+xpc10nz) || (6'd44/*MS*/==-8'd91+xpc10nz) || (6'd44/*MS*/==-8'd90+xpc10nz) || (6'd44/*MS*/==-8'd89+xpc10nz) || (6'd44
              /*MS*/==-8'd88+xpc10nz) || (6'd44/*MS*/==-8'd87+xpc10nz) || (6'd44/*MS*/==-8'd86+xpc10nz) || (6'd44/*MS*/==-8'd85+xpc10nz
              ) || (6'd44/*MS*/==-8'd84+xpc10nz) || (6'd44/*MS*/==-8'd83+xpc10nz) || (6'd44/*MS*/==-8'd82+xpc10nz) || (6'd44/*MS*/==-8'd65
              +xpc10nz) || (6'd44/*MS*/==-8'd64+xpc10nz) || (6'd44/*MS*/==-7'd59+xpc10nz) || (6'd44/*MS*/==-7'd50+xpc10nz) || (6'd44/*MS*/==
              -7'd37+xpc10nz) || (6'd44/*MS*/==-6'd20+xpc10nz) || (6'd44/*MS*/==-6'd19+xpc10nz) || (6'd44/*MS*/==-6'd18+xpc10nz) || (6'd44
              /*MS*/==-6'd17+xpc10nz) || (6'd44/*MS*/==-6'd16+xpc10nz) || (6'd44/*MS*/==-5'd15+xpc10nz) || (6'd44/*MS*/==-5'd14+xpc10nz
              ) || (6'd44/*MS*/==-5'd13+xpc10nz) || (6'd44/*MS*/==-5'd12+xpc10nz) || (6'd44/*MS*/==-5'd11+xpc10nz) || (6'd44/*MS*/==-5'd10
              +xpc10nz) || (6'd44/*MS*/==-5'd9+xpc10nz) || (6'd44/*MS*/==-5'd8+xpc10nz) || (6'd44/*MS*/==-4'd7+xpc10nz) || (6'd44/*MS*/==
              -4'd6+xpc10nz) || (6'd44/*MS*/==-4'd5+xpc10nz) || (6'd44/*MS*/==-4'd4+xpc10nz) || (6'd44/*MS*/==-3'd3+xpc10nz) || (6'd44
              /*MS*/==-3'd2+xpc10nz) || (6'd44/*MS*/==-2'd1+xpc10nz) || (xpc10nz==6'd44/*US*/)) && !xpc10_clear && !xpc10_stall;

               xpc10_trk43 <= ((6'd43/*MS*/==-11'd609+xpc10nz) || (6'd43/*MS*/==-11'd599+xpc10nz) || (6'd43/*MS*/==-11'd588+xpc10nz) || 
              (6'd43/*MS*/==-11'd576+xpc10nz) || (6'd43/*MS*/==-11'd571+xpc10nz) || (6'd43/*MS*/==-11'd565+xpc10nz) || (6'd43/*MS*/==
              -11'd558+xpc10nz) || (6'd43/*MS*/==-11'd550+xpc10nz) || (6'd43/*MS*/==-11'd549+xpc10nz) || (6'd43/*MS*/==-11'd547+xpc10nz
              ) || (6'd43/*MS*/==-11'd544+xpc10nz) || (6'd43/*MS*/==-11'd540+xpc10nz) || (6'd43/*MS*/==-11'd539+xpc10nz) || (6'd43/*MS*/==
              -11'd537+xpc10nz) || (6'd43/*MS*/==-11'd534+xpc10nz) || (6'd43/*MS*/==-11'd532+xpc10nz) || (6'd43/*MS*/==-11'd528+xpc10nz
              ) || (6'd43/*MS*/==-10'd503+xpc10nz) || (6'd43/*MS*/==-10'd502+xpc10nz) || (6'd43/*MS*/==-10'd472+xpc10nz) || (6'd43/*MS*/==
              -10'd407+xpc10nz) || (6'd43/*MS*/==-10'd342+xpc10nz) || (6'd43/*MS*/==-10'd341+xpc10nz) || (6'd43/*MS*/==-10'd340+xpc10nz
              ) || (6'd43/*MS*/==-10'd338+xpc10nz) || (6'd43/*MS*/==-10'd335+xpc10nz) || (6'd43/*MS*/==-10'd334+xpc10nz) || (6'd43/*MS*/==
              -10'd330+xpc10nz) || (6'd43/*MS*/==-10'd329+xpc10nz) || (6'd43/*MS*/==-10'd327+xpc10nz) || (6'd43/*MS*/==-10'd324+xpc10nz
              ) || (6'd43/*MS*/==-10'd323+xpc10nz) || (6'd43/*MS*/==-10'd322+xpc10nz) || (6'd43/*MS*/==-10'd321+xpc10nz) || (6'd43/*MS*/==
              -10'd320+xpc10nz) || (6'd43/*MS*/==-10'd319+xpc10nz) || (6'd43/*MS*/==-10'd318+xpc10nz) || (6'd43/*MS*/==-10'd314+xpc10nz
              ) || (6'd43/*MS*/==-10'd289+xpc10nz) || (6'd43/*MS*/==-10'd287+xpc10nz) || (6'd43/*MS*/==-10'd285+xpc10nz) || (6'd43/*MS*/==
              -10'd284+xpc10nz) || (6'd43/*MS*/==-10'd259+xpc10nz) || (6'd43/*MS*/==-10'd258+xpc10nz) || (6'd43/*MS*/==-10'd257+xpc10nz
              ) || (6'd43/*MS*/==-9'd255+xpc10nz) || (6'd43/*MS*/==-9'd254+xpc10nz) || (6'd43/*MS*/==-9'd253+xpc10nz) || (6'd43/*MS*/==
              -9'd252+xpc10nz) || (6'd43/*MS*/==-9'd251+xpc10nz) || (6'd43/*MS*/==-9'd250+xpc10nz) || (6'd43/*MS*/==-9'd249+xpc10nz) || 
              (6'd43/*MS*/==-9'd248+xpc10nz) || (6'd43/*MS*/==-9'd247+xpc10nz) || (6'd43/*MS*/==-9'd246+xpc10nz) || (6'd43/*MS*/==-9'd245
              +xpc10nz) || (6'd43/*MS*/==-9'd244+xpc10nz) || (6'd43/*MS*/==-9'd242+xpc10nz) || (6'd43/*MS*/==-9'd241+xpc10nz) || (6'd43
              /*MS*/==-9'd239+xpc10nz) || (6'd43/*MS*/==-9'd238+xpc10nz) || (6'd43/*MS*/==-9'd236+xpc10nz) || (6'd43/*MS*/==-9'd171+xpc10nz
              ) || (6'd43/*MS*/==-8'd106+xpc10nz) || (6'd43/*MS*/==-8'd105+xpc10nz) || (6'd43/*MS*/==-8'd104+xpc10nz) || (6'd43/*MS*/==
              -8'd103+xpc10nz) || (6'd43/*MS*/==-8'd102+xpc10nz) || (6'd43/*MS*/==-8'd101+xpc10nz) || (6'd43/*MS*/==-8'd100+xpc10nz) || 
              (6'd43/*MS*/==-8'd99+xpc10nz) || (6'd43/*MS*/==-8'd98+xpc10nz) || (6'd43/*MS*/==-8'd97+xpc10nz) || (6'd43/*MS*/==-8'd96
              +xpc10nz) || (6'd43/*MS*/==-8'd95+xpc10nz) || (6'd43/*MS*/==-8'd94+xpc10nz) || (6'd43/*MS*/==-8'd93+xpc10nz) || (6'd43/*MS*/==
              -8'd92+xpc10nz) || (6'd43/*MS*/==-8'd91+xpc10nz) || (6'd43/*MS*/==-8'd90+xpc10nz) || (6'd43/*MS*/==-8'd89+xpc10nz) || (6'd43
              /*MS*/==-8'd88+xpc10nz) || (6'd43/*MS*/==-8'd87+xpc10nz) || (6'd43/*MS*/==-8'd86+xpc10nz) || (6'd43/*MS*/==-8'd85+xpc10nz
              ) || (6'd43/*MS*/==-8'd84+xpc10nz) || (6'd43/*MS*/==-8'd83+xpc10nz) || (6'd43/*MS*/==-8'd82+xpc10nz) || (6'd43/*MS*/==-8'd65
              +xpc10nz) || (6'd43/*MS*/==-8'd64+xpc10nz) || (6'd43/*MS*/==-7'd59+xpc10nz) || (6'd43/*MS*/==-7'd50+xpc10nz) || (6'd43/*MS*/==
              -7'd37+xpc10nz) || (6'd43/*MS*/==-6'd20+xpc10nz) || (6'd43/*MS*/==-6'd19+xpc10nz) || (6'd43/*MS*/==-6'd18+xpc10nz) || (6'd43
              /*MS*/==-6'd17+xpc10nz) || (6'd43/*MS*/==-6'd16+xpc10nz) || (6'd43/*MS*/==-5'd15+xpc10nz) || (6'd43/*MS*/==-5'd14+xpc10nz
              ) || (6'd43/*MS*/==-5'd13+xpc10nz) || (6'd43/*MS*/==-5'd12+xpc10nz) || (6'd43/*MS*/==-5'd11+xpc10nz) || (6'd43/*MS*/==-5'd10
              +xpc10nz) || (6'd43/*MS*/==-5'd9+xpc10nz) || (6'd43/*MS*/==-5'd8+xpc10nz) || (6'd43/*MS*/==-4'd7+xpc10nz) || (6'd43/*MS*/==
              -4'd6+xpc10nz) || (6'd43/*MS*/==-4'd5+xpc10nz) || (6'd43/*MS*/==-4'd4+xpc10nz) || (6'd43/*MS*/==-3'd3+xpc10nz) || (6'd43
              /*MS*/==-3'd2+xpc10nz) || (6'd43/*MS*/==-2'd1+xpc10nz) || (xpc10nz==6'd43/*US*/)) && !xpc10_clear && !xpc10_stall;

               xpc10_trk42 <= ((6'd42/*MS*/==-11'd609+xpc10nz) || (6'd42/*MS*/==-11'd599+xpc10nz) || (6'd42/*MS*/==-11'd588+xpc10nz) || 
              (6'd42/*MS*/==-11'd576+xpc10nz) || (6'd42/*MS*/==-11'd571+xpc10nz) || (6'd42/*MS*/==-11'd565+xpc10nz) || (6'd42/*MS*/==
              -11'd558+xpc10nz) || (6'd42/*MS*/==-11'd550+xpc10nz) || (6'd42/*MS*/==-11'd549+xpc10nz) || (6'd42/*MS*/==-11'd547+xpc10nz
              ) || (6'd42/*MS*/==-11'd544+xpc10nz) || (6'd42/*MS*/==-11'd540+xpc10nz) || (6'd42/*MS*/==-11'd539+xpc10nz) || (6'd42/*MS*/==
              -11'd537+xpc10nz) || (6'd42/*MS*/==-11'd534+xpc10nz) || (6'd42/*MS*/==-11'd532+xpc10nz) || (6'd42/*MS*/==-11'd528+xpc10nz
              ) || (6'd42/*MS*/==-10'd503+xpc10nz) || (6'd42/*MS*/==-10'd502+xpc10nz) || (6'd42/*MS*/==-10'd472+xpc10nz) || (6'd42/*MS*/==
              -10'd407+xpc10nz) || (6'd42/*MS*/==-10'd342+xpc10nz) || (6'd42/*MS*/==-10'd341+xpc10nz) || (6'd42/*MS*/==-10'd340+xpc10nz
              ) || (6'd42/*MS*/==-10'd338+xpc10nz) || (6'd42/*MS*/==-10'd335+xpc10nz) || (6'd42/*MS*/==-10'd334+xpc10nz) || (6'd42/*MS*/==
              -10'd330+xpc10nz) || (6'd42/*MS*/==-10'd329+xpc10nz) || (6'd42/*MS*/==-10'd327+xpc10nz) || (6'd42/*MS*/==-10'd324+xpc10nz
              ) || (6'd42/*MS*/==-10'd323+xpc10nz) || (6'd42/*MS*/==-10'd322+xpc10nz) || (6'd42/*MS*/==-10'd321+xpc10nz) || (6'd42/*MS*/==
              -10'd320+xpc10nz) || (6'd42/*MS*/==-10'd319+xpc10nz) || (6'd42/*MS*/==-10'd318+xpc10nz) || (6'd42/*MS*/==-10'd314+xpc10nz
              ) || (6'd42/*MS*/==-10'd289+xpc10nz) || (6'd42/*MS*/==-10'd287+xpc10nz) || (6'd42/*MS*/==-10'd285+xpc10nz) || (6'd42/*MS*/==
              -10'd284+xpc10nz) || (6'd42/*MS*/==-10'd259+xpc10nz) || (6'd42/*MS*/==-10'd258+xpc10nz) || (6'd42/*MS*/==-10'd257+xpc10nz
              ) || (6'd42/*MS*/==-9'd255+xpc10nz) || (6'd42/*MS*/==-9'd254+xpc10nz) || (6'd42/*MS*/==-9'd253+xpc10nz) || (6'd42/*MS*/==
              -9'd252+xpc10nz) || (6'd42/*MS*/==-9'd251+xpc10nz) || (6'd42/*MS*/==-9'd250+xpc10nz) || (6'd42/*MS*/==-9'd249+xpc10nz) || 
              (6'd42/*MS*/==-9'd248+xpc10nz) || (6'd42/*MS*/==-9'd247+xpc10nz) || (6'd42/*MS*/==-9'd246+xpc10nz) || (6'd42/*MS*/==-9'd245
              +xpc10nz) || (6'd42/*MS*/==-9'd244+xpc10nz) || (6'd42/*MS*/==-9'd242+xpc10nz) || (6'd42/*MS*/==-9'd241+xpc10nz) || (6'd42
              /*MS*/==-9'd239+xpc10nz) || (6'd42/*MS*/==-9'd238+xpc10nz) || (6'd42/*MS*/==-9'd236+xpc10nz) || (6'd42/*MS*/==-9'd171+xpc10nz
              ) || (6'd42/*MS*/==-8'd106+xpc10nz) || (6'd42/*MS*/==-8'd105+xpc10nz) || (6'd42/*MS*/==-8'd104+xpc10nz) || (6'd42/*MS*/==
              -8'd103+xpc10nz) || (6'd42/*MS*/==-8'd102+xpc10nz) || (6'd42/*MS*/==-8'd101+xpc10nz) || (6'd42/*MS*/==-8'd100+xpc10nz) || 
              (6'd42/*MS*/==-8'd99+xpc10nz) || (6'd42/*MS*/==-8'd98+xpc10nz) || (6'd42/*MS*/==-8'd97+xpc10nz) || (6'd42/*MS*/==-8'd96
              +xpc10nz) || (6'd42/*MS*/==-8'd95+xpc10nz) || (6'd42/*MS*/==-8'd94+xpc10nz) || (6'd42/*MS*/==-8'd93+xpc10nz) || (6'd42/*MS*/==
              -8'd92+xpc10nz) || (6'd42/*MS*/==-8'd91+xpc10nz) || (6'd42/*MS*/==-8'd90+xpc10nz) || (6'd42/*MS*/==-8'd89+xpc10nz) || (6'd42
              /*MS*/==-8'd88+xpc10nz) || (6'd42/*MS*/==-8'd87+xpc10nz) || (6'd42/*MS*/==-8'd86+xpc10nz) || (6'd42/*MS*/==-8'd85+xpc10nz
              ) || (6'd42/*MS*/==-8'd84+xpc10nz) || (6'd42/*MS*/==-8'd83+xpc10nz) || (6'd42/*MS*/==-8'd82+xpc10nz) || (6'd42/*MS*/==-8'd65
              +xpc10nz) || (6'd42/*MS*/==-8'd64+xpc10nz) || (6'd42/*MS*/==-7'd59+xpc10nz) || (6'd42/*MS*/==-7'd50+xpc10nz) || (6'd42/*MS*/==
              -7'd37+xpc10nz) || (6'd42/*MS*/==-6'd20+xpc10nz) || (6'd42/*MS*/==-6'd19+xpc10nz) || (6'd42/*MS*/==-6'd18+xpc10nz) || (6'd42
              /*MS*/==-6'd17+xpc10nz) || (6'd42/*MS*/==-6'd16+xpc10nz) || (6'd42/*MS*/==-5'd15+xpc10nz) || (6'd42/*MS*/==-5'd14+xpc10nz
              ) || (6'd42/*MS*/==-5'd13+xpc10nz) || (6'd42/*MS*/==-5'd12+xpc10nz) || (6'd42/*MS*/==-5'd11+xpc10nz) || (6'd42/*MS*/==-5'd10
              +xpc10nz) || (6'd42/*MS*/==-5'd9+xpc10nz) || (6'd42/*MS*/==-5'd8+xpc10nz) || (6'd42/*MS*/==-4'd7+xpc10nz) || (6'd42/*MS*/==
              -4'd6+xpc10nz) || (6'd42/*MS*/==-4'd5+xpc10nz) || (6'd42/*MS*/==-4'd4+xpc10nz) || (6'd42/*MS*/==-3'd3+xpc10nz) || (6'd42
              /*MS*/==-3'd2+xpc10nz) || (6'd42/*MS*/==-2'd1+xpc10nz) || (xpc10nz==6'd42/*US*/)) && !xpc10_clear && !xpc10_stall;

               xpc10_trk41 <= ((6'd41/*MS*/==-11'd609+xpc10nz) || (6'd41/*MS*/==-11'd599+xpc10nz) || (6'd41/*MS*/==-11'd588+xpc10nz) || 
              (6'd41/*MS*/==-11'd576+xpc10nz) || (6'd41/*MS*/==-11'd571+xpc10nz) || (6'd41/*MS*/==-11'd565+xpc10nz) || (6'd41/*MS*/==
              -11'd558+xpc10nz) || (6'd41/*MS*/==-11'd550+xpc10nz) || (6'd41/*MS*/==-11'd549+xpc10nz) || (6'd41/*MS*/==-11'd547+xpc10nz
              ) || (6'd41/*MS*/==-11'd544+xpc10nz) || (6'd41/*MS*/==-11'd540+xpc10nz) || (6'd41/*MS*/==-11'd539+xpc10nz) || (6'd41/*MS*/==
              -11'd537+xpc10nz) || (6'd41/*MS*/==-11'd534+xpc10nz) || (6'd41/*MS*/==-11'd532+xpc10nz) || (6'd41/*MS*/==-11'd528+xpc10nz
              ) || (6'd41/*MS*/==-10'd503+xpc10nz) || (6'd41/*MS*/==-10'd502+xpc10nz) || (6'd41/*MS*/==-10'd472+xpc10nz) || (6'd41/*MS*/==
              -10'd407+xpc10nz) || (6'd41/*MS*/==-10'd342+xpc10nz) || (6'd41/*MS*/==-10'd341+xpc10nz) || (6'd41/*MS*/==-10'd340+xpc10nz
              ) || (6'd41/*MS*/==-10'd338+xpc10nz) || (6'd41/*MS*/==-10'd335+xpc10nz) || (6'd41/*MS*/==-10'd334+xpc10nz) || (6'd41/*MS*/==
              -10'd330+xpc10nz) || (6'd41/*MS*/==-10'd329+xpc10nz) || (6'd41/*MS*/==-10'd327+xpc10nz) || (6'd41/*MS*/==-10'd324+xpc10nz
              ) || (6'd41/*MS*/==-10'd323+xpc10nz) || (6'd41/*MS*/==-10'd322+xpc10nz) || (6'd41/*MS*/==-10'd321+xpc10nz) || (6'd41/*MS*/==
              -10'd320+xpc10nz) || (6'd41/*MS*/==-10'd319+xpc10nz) || (6'd41/*MS*/==-10'd318+xpc10nz) || (6'd41/*MS*/==-10'd314+xpc10nz
              ) || (6'd41/*MS*/==-10'd289+xpc10nz) || (6'd41/*MS*/==-10'd287+xpc10nz) || (6'd41/*MS*/==-10'd285+xpc10nz) || (6'd41/*MS*/==
              -10'd284+xpc10nz) || (6'd41/*MS*/==-10'd259+xpc10nz) || (6'd41/*MS*/==-10'd258+xpc10nz) || (6'd41/*MS*/==-10'd257+xpc10nz
              ) || (6'd41/*MS*/==-9'd255+xpc10nz) || (6'd41/*MS*/==-9'd254+xpc10nz) || (6'd41/*MS*/==-9'd253+xpc10nz) || (6'd41/*MS*/==
              -9'd252+xpc10nz) || (6'd41/*MS*/==-9'd251+xpc10nz) || (6'd41/*MS*/==-9'd250+xpc10nz) || (6'd41/*MS*/==-9'd249+xpc10nz) || 
              (6'd41/*MS*/==-9'd248+xpc10nz) || (6'd41/*MS*/==-9'd247+xpc10nz) || (6'd41/*MS*/==-9'd246+xpc10nz) || (6'd41/*MS*/==-9'd245
              +xpc10nz) || (6'd41/*MS*/==-9'd244+xpc10nz) || (6'd41/*MS*/==-9'd242+xpc10nz) || (6'd41/*MS*/==-9'd241+xpc10nz) || (6'd41
              /*MS*/==-9'd239+xpc10nz) || (6'd41/*MS*/==-9'd238+xpc10nz) || (6'd41/*MS*/==-9'd236+xpc10nz) || (6'd41/*MS*/==-9'd171+xpc10nz
              ) || (6'd41/*MS*/==-8'd106+xpc10nz) || (6'd41/*MS*/==-8'd105+xpc10nz) || (6'd41/*MS*/==-8'd104+xpc10nz) || (6'd41/*MS*/==
              -8'd103+xpc10nz) || (6'd41/*MS*/==-8'd102+xpc10nz) || (6'd41/*MS*/==-8'd101+xpc10nz) || (6'd41/*MS*/==-8'd100+xpc10nz) || 
              (6'd41/*MS*/==-8'd99+xpc10nz) || (6'd41/*MS*/==-8'd98+xpc10nz) || (6'd41/*MS*/==-8'd97+xpc10nz) || (6'd41/*MS*/==-8'd96
              +xpc10nz) || (6'd41/*MS*/==-8'd95+xpc10nz) || (6'd41/*MS*/==-8'd94+xpc10nz) || (6'd41/*MS*/==-8'd93+xpc10nz) || (6'd41/*MS*/==
              -8'd92+xpc10nz) || (6'd41/*MS*/==-8'd91+xpc10nz) || (6'd41/*MS*/==-8'd90+xpc10nz) || (6'd41/*MS*/==-8'd89+xpc10nz) || (6'd41
              /*MS*/==-8'd88+xpc10nz) || (6'd41/*MS*/==-8'd87+xpc10nz) || (6'd41/*MS*/==-8'd86+xpc10nz) || (6'd41/*MS*/==-8'd85+xpc10nz
              ) || (6'd41/*MS*/==-8'd84+xpc10nz) || (6'd41/*MS*/==-8'd83+xpc10nz) || (6'd41/*MS*/==-8'd82+xpc10nz) || (6'd41/*MS*/==-8'd65
              +xpc10nz) || (6'd41/*MS*/==-8'd64+xpc10nz) || (6'd41/*MS*/==-7'd59+xpc10nz) || (6'd41/*MS*/==-7'd50+xpc10nz) || (6'd41/*MS*/==
              -7'd37+xpc10nz) || (6'd41/*MS*/==-6'd20+xpc10nz) || (6'd41/*MS*/==-6'd19+xpc10nz) || (6'd41/*MS*/==-6'd18+xpc10nz) || (6'd41
              /*MS*/==-6'd17+xpc10nz) || (6'd41/*MS*/==-6'd16+xpc10nz) || (6'd41/*MS*/==-5'd15+xpc10nz) || (6'd41/*MS*/==-5'd14+xpc10nz
              ) || (6'd41/*MS*/==-5'd13+xpc10nz) || (6'd41/*MS*/==-5'd12+xpc10nz) || (6'd41/*MS*/==-5'd11+xpc10nz) || (6'd41/*MS*/==-5'd10
              +xpc10nz) || (6'd41/*MS*/==-5'd9+xpc10nz) || (6'd41/*MS*/==-5'd8+xpc10nz) || (6'd41/*MS*/==-4'd7+xpc10nz) || (6'd41/*MS*/==
              -4'd6+xpc10nz) || (6'd41/*MS*/==-4'd5+xpc10nz) || (6'd41/*MS*/==-4'd4+xpc10nz) || (6'd41/*MS*/==-3'd3+xpc10nz) || (6'd41
              /*MS*/==-3'd2+xpc10nz) || (6'd41/*MS*/==-2'd1+xpc10nz) || (xpc10nz==6'd41/*US*/)) && !xpc10_clear && !xpc10_stall;

               xpc10_trk40 <= ((6'd40/*MS*/==-11'd609+xpc10nz) || (6'd40/*MS*/==-11'd599+xpc10nz) || (6'd40/*MS*/==-11'd588+xpc10nz) || 
              (6'd40/*MS*/==-11'd576+xpc10nz) || (6'd40/*MS*/==-11'd571+xpc10nz) || (6'd40/*MS*/==-11'd565+xpc10nz) || (6'd40/*MS*/==
              -11'd558+xpc10nz) || (6'd40/*MS*/==-11'd550+xpc10nz) || (6'd40/*MS*/==-11'd549+xpc10nz) || (6'd40/*MS*/==-11'd547+xpc10nz
              ) || (6'd40/*MS*/==-11'd544+xpc10nz) || (6'd40/*MS*/==-11'd540+xpc10nz) || (6'd40/*MS*/==-11'd539+xpc10nz) || (6'd40/*MS*/==
              -11'd537+xpc10nz) || (6'd40/*MS*/==-11'd534+xpc10nz) || (6'd40/*MS*/==-11'd532+xpc10nz) || (6'd40/*MS*/==-11'd528+xpc10nz
              ) || (6'd40/*MS*/==-10'd503+xpc10nz) || (6'd40/*MS*/==-10'd502+xpc10nz) || (6'd40/*MS*/==-10'd472+xpc10nz) || (6'd40/*MS*/==
              -10'd407+xpc10nz) || (6'd40/*MS*/==-10'd342+xpc10nz) || (6'd40/*MS*/==-10'd341+xpc10nz) || (6'd40/*MS*/==-10'd340+xpc10nz
              ) || (6'd40/*MS*/==-10'd338+xpc10nz) || (6'd40/*MS*/==-10'd335+xpc10nz) || (6'd40/*MS*/==-10'd334+xpc10nz) || (6'd40/*MS*/==
              -10'd330+xpc10nz) || (6'd40/*MS*/==-10'd329+xpc10nz) || (6'd40/*MS*/==-10'd327+xpc10nz) || (6'd40/*MS*/==-10'd324+xpc10nz
              ) || (6'd40/*MS*/==-10'd323+xpc10nz) || (6'd40/*MS*/==-10'd322+xpc10nz) || (6'd40/*MS*/==-10'd321+xpc10nz) || (6'd40/*MS*/==
              -10'd320+xpc10nz) || (6'd40/*MS*/==-10'd319+xpc10nz) || (6'd40/*MS*/==-10'd318+xpc10nz) || (6'd40/*MS*/==-10'd314+xpc10nz
              ) || (6'd40/*MS*/==-10'd289+xpc10nz) || (6'd40/*MS*/==-10'd287+xpc10nz) || (6'd40/*MS*/==-10'd285+xpc10nz) || (6'd40/*MS*/==
              -10'd284+xpc10nz) || (6'd40/*MS*/==-10'd259+xpc10nz) || (6'd40/*MS*/==-10'd258+xpc10nz) || (6'd40/*MS*/==-10'd257+xpc10nz
              ) || (6'd40/*MS*/==-9'd255+xpc10nz) || (6'd40/*MS*/==-9'd254+xpc10nz) || (6'd40/*MS*/==-9'd253+xpc10nz) || (6'd40/*MS*/==
              -9'd252+xpc10nz) || (6'd40/*MS*/==-9'd251+xpc10nz) || (6'd40/*MS*/==-9'd250+xpc10nz) || (6'd40/*MS*/==-9'd249+xpc10nz) || 
              (6'd40/*MS*/==-9'd248+xpc10nz) || (6'd40/*MS*/==-9'd247+xpc10nz) || (6'd40/*MS*/==-9'd246+xpc10nz) || (6'd40/*MS*/==-9'd245
              +xpc10nz) || (6'd40/*MS*/==-9'd244+xpc10nz) || (6'd40/*MS*/==-9'd242+xpc10nz) || (6'd40/*MS*/==-9'd241+xpc10nz) || (6'd40
              /*MS*/==-9'd239+xpc10nz) || (6'd40/*MS*/==-9'd238+xpc10nz) || (6'd40/*MS*/==-9'd236+xpc10nz) || (6'd40/*MS*/==-9'd171+xpc10nz
              ) || (6'd40/*MS*/==-8'd106+xpc10nz) || (6'd40/*MS*/==-8'd105+xpc10nz) || (6'd40/*MS*/==-8'd104+xpc10nz) || (6'd40/*MS*/==
              -8'd103+xpc10nz) || (6'd40/*MS*/==-8'd102+xpc10nz) || (6'd40/*MS*/==-8'd101+xpc10nz) || (6'd40/*MS*/==-8'd100+xpc10nz) || 
              (6'd40/*MS*/==-8'd99+xpc10nz) || (6'd40/*MS*/==-8'd98+xpc10nz) || (6'd40/*MS*/==-8'd97+xpc10nz) || (6'd40/*MS*/==-8'd96
              +xpc10nz) || (6'd40/*MS*/==-8'd95+xpc10nz) || (6'd40/*MS*/==-8'd94+xpc10nz) || (6'd40/*MS*/==-8'd93+xpc10nz) || (6'd40/*MS*/==
              -8'd92+xpc10nz) || (6'd40/*MS*/==-8'd91+xpc10nz) || (6'd40/*MS*/==-8'd90+xpc10nz) || (6'd40/*MS*/==-8'd89+xpc10nz) || (6'd40
              /*MS*/==-8'd88+xpc10nz) || (6'd40/*MS*/==-8'd87+xpc10nz) || (6'd40/*MS*/==-8'd86+xpc10nz) || (6'd40/*MS*/==-8'd85+xpc10nz
              ) || (6'd40/*MS*/==-8'd84+xpc10nz) || (6'd40/*MS*/==-8'd83+xpc10nz) || (6'd40/*MS*/==-8'd82+xpc10nz) || (6'd40/*MS*/==-8'd65
              +xpc10nz) || (6'd40/*MS*/==-8'd64+xpc10nz) || (6'd40/*MS*/==-7'd59+xpc10nz) || (6'd40/*MS*/==-7'd50+xpc10nz) || (6'd40/*MS*/==
              -7'd37+xpc10nz) || (6'd40/*MS*/==-6'd20+xpc10nz) || (6'd40/*MS*/==-6'd19+xpc10nz) || (6'd40/*MS*/==-6'd18+xpc10nz) || (6'd40
              /*MS*/==-6'd17+xpc10nz) || (6'd40/*MS*/==-6'd16+xpc10nz) || (6'd40/*MS*/==-5'd15+xpc10nz) || (6'd40/*MS*/==-5'd14+xpc10nz
              ) || (6'd40/*MS*/==-5'd13+xpc10nz) || (6'd40/*MS*/==-5'd12+xpc10nz) || (6'd40/*MS*/==-5'd11+xpc10nz) || (6'd40/*MS*/==-5'd10
              +xpc10nz) || (6'd40/*MS*/==-5'd9+xpc10nz) || (6'd40/*MS*/==-5'd8+xpc10nz) || (6'd40/*MS*/==-4'd7+xpc10nz) || (6'd40/*MS*/==
              -4'd6+xpc10nz) || (6'd40/*MS*/==-4'd5+xpc10nz) || (6'd40/*MS*/==-4'd4+xpc10nz) || (6'd40/*MS*/==-3'd3+xpc10nz) || (6'd40
              /*MS*/==-3'd2+xpc10nz) || (6'd40/*MS*/==-2'd1+xpc10nz) || (xpc10nz==6'd40/*US*/)) && !xpc10_clear && !xpc10_stall;

               xpc10_trk39 <= ((6'd39/*MS*/==-11'd609+xpc10nz) || (6'd39/*MS*/==-11'd599+xpc10nz) || (6'd39/*MS*/==-11'd588+xpc10nz) || 
              (6'd39/*MS*/==-11'd576+xpc10nz) || (6'd39/*MS*/==-11'd571+xpc10nz) || (6'd39/*MS*/==-11'd565+xpc10nz) || (6'd39/*MS*/==
              -11'd558+xpc10nz) || (6'd39/*MS*/==-11'd550+xpc10nz) || (6'd39/*MS*/==-11'd549+xpc10nz) || (6'd39/*MS*/==-11'd547+xpc10nz
              ) || (6'd39/*MS*/==-11'd544+xpc10nz) || (6'd39/*MS*/==-11'd540+xpc10nz) || (6'd39/*MS*/==-11'd539+xpc10nz) || (6'd39/*MS*/==
              -11'd537+xpc10nz) || (6'd39/*MS*/==-11'd534+xpc10nz) || (6'd39/*MS*/==-11'd532+xpc10nz) || (6'd39/*MS*/==-11'd528+xpc10nz
              ) || (6'd39/*MS*/==-10'd503+xpc10nz) || (6'd39/*MS*/==-10'd502+xpc10nz) || (6'd39/*MS*/==-10'd472+xpc10nz) || (6'd39/*MS*/==
              -10'd407+xpc10nz) || (6'd39/*MS*/==-10'd342+xpc10nz) || (6'd39/*MS*/==-10'd341+xpc10nz) || (6'd39/*MS*/==-10'd340+xpc10nz
              ) || (6'd39/*MS*/==-10'd338+xpc10nz) || (6'd39/*MS*/==-10'd335+xpc10nz) || (6'd39/*MS*/==-10'd334+xpc10nz) || (6'd39/*MS*/==
              -10'd330+xpc10nz) || (6'd39/*MS*/==-10'd329+xpc10nz) || (6'd39/*MS*/==-10'd327+xpc10nz) || (6'd39/*MS*/==-10'd324+xpc10nz
              ) || (6'd39/*MS*/==-10'd323+xpc10nz) || (6'd39/*MS*/==-10'd322+xpc10nz) || (6'd39/*MS*/==-10'd321+xpc10nz) || (6'd39/*MS*/==
              -10'd320+xpc10nz) || (6'd39/*MS*/==-10'd319+xpc10nz) || (6'd39/*MS*/==-10'd318+xpc10nz) || (6'd39/*MS*/==-10'd314+xpc10nz
              ) || (6'd39/*MS*/==-10'd289+xpc10nz) || (6'd39/*MS*/==-10'd287+xpc10nz) || (6'd39/*MS*/==-10'd285+xpc10nz) || (6'd39/*MS*/==
              -10'd284+xpc10nz) || (6'd39/*MS*/==-10'd259+xpc10nz) || (6'd39/*MS*/==-10'd258+xpc10nz) || (6'd39/*MS*/==-10'd257+xpc10nz
              ) || (6'd39/*MS*/==-9'd255+xpc10nz) || (6'd39/*MS*/==-9'd254+xpc10nz) || (6'd39/*MS*/==-9'd253+xpc10nz) || (6'd39/*MS*/==
              -9'd252+xpc10nz) || (6'd39/*MS*/==-9'd251+xpc10nz) || (6'd39/*MS*/==-9'd250+xpc10nz) || (6'd39/*MS*/==-9'd249+xpc10nz) || 
              (6'd39/*MS*/==-9'd248+xpc10nz) || (6'd39/*MS*/==-9'd247+xpc10nz) || (6'd39/*MS*/==-9'd246+xpc10nz) || (6'd39/*MS*/==-9'd245
              +xpc10nz) || (6'd39/*MS*/==-9'd244+xpc10nz) || (6'd39/*MS*/==-9'd242+xpc10nz) || (6'd39/*MS*/==-9'd241+xpc10nz) || (6'd39
              /*MS*/==-9'd239+xpc10nz) || (6'd39/*MS*/==-9'd238+xpc10nz) || (6'd39/*MS*/==-9'd236+xpc10nz) || (6'd39/*MS*/==-9'd171+xpc10nz
              ) || (6'd39/*MS*/==-8'd106+xpc10nz) || (6'd39/*MS*/==-8'd105+xpc10nz) || (6'd39/*MS*/==-8'd104+xpc10nz) || (6'd39/*MS*/==
              -8'd103+xpc10nz) || (6'd39/*MS*/==-8'd102+xpc10nz) || (6'd39/*MS*/==-8'd101+xpc10nz) || (6'd39/*MS*/==-8'd100+xpc10nz) || 
              (6'd39/*MS*/==-8'd99+xpc10nz) || (6'd39/*MS*/==-8'd98+xpc10nz) || (6'd39/*MS*/==-8'd97+xpc10nz) || (6'd39/*MS*/==-8'd96
              +xpc10nz) || (6'd39/*MS*/==-8'd95+xpc10nz) || (6'd39/*MS*/==-8'd94+xpc10nz) || (6'd39/*MS*/==-8'd93+xpc10nz) || (6'd39/*MS*/==
              -8'd92+xpc10nz) || (6'd39/*MS*/==-8'd91+xpc10nz) || (6'd39/*MS*/==-8'd90+xpc10nz) || (6'd39/*MS*/==-8'd89+xpc10nz) || (6'd39
              /*MS*/==-8'd88+xpc10nz) || (6'd39/*MS*/==-8'd87+xpc10nz) || (6'd39/*MS*/==-8'd86+xpc10nz) || (6'd39/*MS*/==-8'd85+xpc10nz
              ) || (6'd39/*MS*/==-8'd84+xpc10nz) || (6'd39/*MS*/==-8'd83+xpc10nz) || (6'd39/*MS*/==-8'd82+xpc10nz) || (6'd39/*MS*/==-8'd65
              +xpc10nz) || (6'd39/*MS*/==-8'd64+xpc10nz) || (6'd39/*MS*/==-7'd59+xpc10nz) || (6'd39/*MS*/==-7'd50+xpc10nz) || (6'd39/*MS*/==
              -7'd37+xpc10nz) || (6'd39/*MS*/==-6'd20+xpc10nz) || (6'd39/*MS*/==-6'd19+xpc10nz) || (6'd39/*MS*/==-6'd18+xpc10nz) || (6'd39
              /*MS*/==-6'd17+xpc10nz) || (6'd39/*MS*/==-6'd16+xpc10nz) || (6'd39/*MS*/==-5'd15+xpc10nz) || (6'd39/*MS*/==-5'd14+xpc10nz
              ) || (6'd39/*MS*/==-5'd13+xpc10nz) || (6'd39/*MS*/==-5'd12+xpc10nz) || (6'd39/*MS*/==-5'd11+xpc10nz) || (6'd39/*MS*/==-5'd10
              +xpc10nz) || (6'd39/*MS*/==-5'd9+xpc10nz) || (6'd39/*MS*/==-5'd8+xpc10nz) || (6'd39/*MS*/==-4'd7+xpc10nz) || (6'd39/*MS*/==
              -4'd6+xpc10nz) || (6'd39/*MS*/==-4'd5+xpc10nz) || (6'd39/*MS*/==-4'd4+xpc10nz) || (6'd39/*MS*/==-3'd3+xpc10nz) || (6'd39
              /*MS*/==-3'd2+xpc10nz) || (6'd39/*MS*/==-2'd1+xpc10nz) || (xpc10nz==6'd39/*US*/)) && !xpc10_clear && !xpc10_stall;

               xpc10_trk38 <= ((6'd38/*MS*/==-11'd609+xpc10nz) || (6'd38/*MS*/==-11'd599+xpc10nz) || (6'd38/*MS*/==-11'd588+xpc10nz) || 
              (6'd38/*MS*/==-11'd576+xpc10nz) || (6'd38/*MS*/==-11'd571+xpc10nz) || (6'd38/*MS*/==-11'd565+xpc10nz) || (6'd38/*MS*/==
              -11'd558+xpc10nz) || (6'd38/*MS*/==-11'd550+xpc10nz) || (6'd38/*MS*/==-11'd549+xpc10nz) || (6'd38/*MS*/==-11'd547+xpc10nz
              ) || (6'd38/*MS*/==-11'd544+xpc10nz) || (6'd38/*MS*/==-11'd540+xpc10nz) || (6'd38/*MS*/==-11'd539+xpc10nz) || (6'd38/*MS*/==
              -11'd537+xpc10nz) || (6'd38/*MS*/==-11'd534+xpc10nz) || (6'd38/*MS*/==-11'd532+xpc10nz) || (6'd38/*MS*/==-11'd528+xpc10nz
              ) || (6'd38/*MS*/==-10'd503+xpc10nz) || (6'd38/*MS*/==-10'd502+xpc10nz) || (6'd38/*MS*/==-10'd472+xpc10nz) || (6'd38/*MS*/==
              -10'd407+xpc10nz) || (6'd38/*MS*/==-10'd342+xpc10nz) || (6'd38/*MS*/==-10'd341+xpc10nz) || (6'd38/*MS*/==-10'd340+xpc10nz
              ) || (6'd38/*MS*/==-10'd338+xpc10nz) || (6'd38/*MS*/==-10'd335+xpc10nz) || (6'd38/*MS*/==-10'd334+xpc10nz) || (6'd38/*MS*/==
              -10'd330+xpc10nz) || (6'd38/*MS*/==-10'd329+xpc10nz) || (6'd38/*MS*/==-10'd327+xpc10nz) || (6'd38/*MS*/==-10'd324+xpc10nz
              ) || (6'd38/*MS*/==-10'd323+xpc10nz) || (6'd38/*MS*/==-10'd322+xpc10nz) || (6'd38/*MS*/==-10'd321+xpc10nz) || (6'd38/*MS*/==
              -10'd320+xpc10nz) || (6'd38/*MS*/==-10'd319+xpc10nz) || (6'd38/*MS*/==-10'd318+xpc10nz) || (6'd38/*MS*/==-10'd314+xpc10nz
              ) || (6'd38/*MS*/==-10'd289+xpc10nz) || (6'd38/*MS*/==-10'd287+xpc10nz) || (6'd38/*MS*/==-10'd285+xpc10nz) || (6'd38/*MS*/==
              -10'd284+xpc10nz) || (6'd38/*MS*/==-10'd259+xpc10nz) || (6'd38/*MS*/==-10'd258+xpc10nz) || (6'd38/*MS*/==-10'd257+xpc10nz
              ) || (6'd38/*MS*/==-9'd255+xpc10nz) || (6'd38/*MS*/==-9'd254+xpc10nz) || (6'd38/*MS*/==-9'd253+xpc10nz) || (6'd38/*MS*/==
              -9'd252+xpc10nz) || (6'd38/*MS*/==-9'd251+xpc10nz) || (6'd38/*MS*/==-9'd250+xpc10nz) || (6'd38/*MS*/==-9'd249+xpc10nz) || 
              (6'd38/*MS*/==-9'd248+xpc10nz) || (6'd38/*MS*/==-9'd247+xpc10nz) || (6'd38/*MS*/==-9'd246+xpc10nz) || (6'd38/*MS*/==-9'd245
              +xpc10nz) || (6'd38/*MS*/==-9'd244+xpc10nz) || (6'd38/*MS*/==-9'd242+xpc10nz) || (6'd38/*MS*/==-9'd241+xpc10nz) || (6'd38
              /*MS*/==-9'd239+xpc10nz) || (6'd38/*MS*/==-9'd238+xpc10nz) || (6'd38/*MS*/==-9'd236+xpc10nz) || (6'd38/*MS*/==-9'd171+xpc10nz
              ) || (6'd38/*MS*/==-8'd106+xpc10nz) || (6'd38/*MS*/==-8'd105+xpc10nz) || (6'd38/*MS*/==-8'd104+xpc10nz) || (6'd38/*MS*/==
              -8'd103+xpc10nz) || (6'd38/*MS*/==-8'd102+xpc10nz) || (6'd38/*MS*/==-8'd101+xpc10nz) || (6'd38/*MS*/==-8'd100+xpc10nz) || 
              (6'd38/*MS*/==-8'd99+xpc10nz) || (6'd38/*MS*/==-8'd98+xpc10nz) || (6'd38/*MS*/==-8'd97+xpc10nz) || (6'd38/*MS*/==-8'd96
              +xpc10nz) || (6'd38/*MS*/==-8'd95+xpc10nz) || (6'd38/*MS*/==-8'd94+xpc10nz) || (6'd38/*MS*/==-8'd93+xpc10nz) || (6'd38/*MS*/==
              -8'd92+xpc10nz) || (6'd38/*MS*/==-8'd91+xpc10nz) || (6'd38/*MS*/==-8'd90+xpc10nz) || (6'd38/*MS*/==-8'd89+xpc10nz) || (6'd38
              /*MS*/==-8'd88+xpc10nz) || (6'd38/*MS*/==-8'd87+xpc10nz) || (6'd38/*MS*/==-8'd86+xpc10nz) || (6'd38/*MS*/==-8'd85+xpc10nz
              ) || (6'd38/*MS*/==-8'd84+xpc10nz) || (6'd38/*MS*/==-8'd83+xpc10nz) || (6'd38/*MS*/==-8'd82+xpc10nz) || (6'd38/*MS*/==-8'd65
              +xpc10nz) || (6'd38/*MS*/==-8'd64+xpc10nz) || (6'd38/*MS*/==-7'd59+xpc10nz) || (6'd38/*MS*/==-7'd50+xpc10nz) || (6'd38/*MS*/==
              -7'd37+xpc10nz) || (6'd38/*MS*/==-6'd20+xpc10nz) || (6'd38/*MS*/==-6'd19+xpc10nz) || (6'd38/*MS*/==-6'd18+xpc10nz) || (6'd38
              /*MS*/==-6'd17+xpc10nz) || (6'd38/*MS*/==-6'd16+xpc10nz) || (6'd38/*MS*/==-5'd15+xpc10nz) || (6'd38/*MS*/==-5'd14+xpc10nz
              ) || (6'd38/*MS*/==-5'd13+xpc10nz) || (6'd38/*MS*/==-5'd12+xpc10nz) || (6'd38/*MS*/==-5'd11+xpc10nz) || (6'd38/*MS*/==-5'd10
              +xpc10nz) || (6'd38/*MS*/==-5'd9+xpc10nz) || (6'd38/*MS*/==-5'd8+xpc10nz) || (6'd38/*MS*/==-4'd7+xpc10nz) || (6'd38/*MS*/==
              -4'd6+xpc10nz) || (6'd38/*MS*/==-4'd5+xpc10nz) || (6'd38/*MS*/==-4'd4+xpc10nz) || (6'd38/*MS*/==-3'd3+xpc10nz) || (6'd38
              /*MS*/==-3'd2+xpc10nz) || (6'd38/*MS*/==-2'd1+xpc10nz) || (xpc10nz==6'd38/*US*/)) && !xpc10_clear && !xpc10_stall;

               xpc10_trk37 <= ((6'd37/*MS*/==-11'd609+xpc10nz) || (6'd37/*MS*/==-11'd599+xpc10nz) || (6'd37/*MS*/==-11'd588+xpc10nz) || 
              (6'd37/*MS*/==-11'd576+xpc10nz) || (6'd37/*MS*/==-11'd571+xpc10nz) || (6'd37/*MS*/==-11'd565+xpc10nz) || (6'd37/*MS*/==
              -11'd558+xpc10nz) || (6'd37/*MS*/==-11'd550+xpc10nz) || (6'd37/*MS*/==-11'd549+xpc10nz) || (6'd37/*MS*/==-11'd547+xpc10nz
              ) || (6'd37/*MS*/==-11'd544+xpc10nz) || (6'd37/*MS*/==-11'd540+xpc10nz) || (6'd37/*MS*/==-11'd539+xpc10nz) || (6'd37/*MS*/==
              -11'd537+xpc10nz) || (6'd37/*MS*/==-11'd534+xpc10nz) || (6'd37/*MS*/==-11'd532+xpc10nz) || (6'd37/*MS*/==-11'd528+xpc10nz
              ) || (6'd37/*MS*/==-10'd503+xpc10nz) || (6'd37/*MS*/==-10'd502+xpc10nz) || (6'd37/*MS*/==-10'd472+xpc10nz) || (6'd37/*MS*/==
              -10'd407+xpc10nz) || (6'd37/*MS*/==-10'd342+xpc10nz) || (6'd37/*MS*/==-10'd341+xpc10nz) || (6'd37/*MS*/==-10'd340+xpc10nz
              ) || (6'd37/*MS*/==-10'd338+xpc10nz) || (6'd37/*MS*/==-10'd335+xpc10nz) || (6'd37/*MS*/==-10'd334+xpc10nz) || (6'd37/*MS*/==
              -10'd330+xpc10nz) || (6'd37/*MS*/==-10'd329+xpc10nz) || (6'd37/*MS*/==-10'd327+xpc10nz) || (6'd37/*MS*/==-10'd324+xpc10nz
              ) || (6'd37/*MS*/==-10'd323+xpc10nz) || (6'd37/*MS*/==-10'd322+xpc10nz) || (6'd37/*MS*/==-10'd321+xpc10nz) || (6'd37/*MS*/==
              -10'd320+xpc10nz) || (6'd37/*MS*/==-10'd319+xpc10nz) || (6'd37/*MS*/==-10'd318+xpc10nz) || (6'd37/*MS*/==-10'd314+xpc10nz
              ) || (6'd37/*MS*/==-10'd289+xpc10nz) || (6'd37/*MS*/==-10'd287+xpc10nz) || (6'd37/*MS*/==-10'd285+xpc10nz) || (6'd37/*MS*/==
              -10'd284+xpc10nz) || (6'd37/*MS*/==-10'd259+xpc10nz) || (6'd37/*MS*/==-10'd258+xpc10nz) || (6'd37/*MS*/==-10'd257+xpc10nz
              ) || (6'd37/*MS*/==-9'd255+xpc10nz) || (6'd37/*MS*/==-9'd254+xpc10nz) || (6'd37/*MS*/==-9'd253+xpc10nz) || (6'd37/*MS*/==
              -9'd252+xpc10nz) || (6'd37/*MS*/==-9'd251+xpc10nz) || (6'd37/*MS*/==-9'd250+xpc10nz) || (6'd37/*MS*/==-9'd249+xpc10nz) || 
              (6'd37/*MS*/==-9'd248+xpc10nz) || (6'd37/*MS*/==-9'd247+xpc10nz) || (6'd37/*MS*/==-9'd246+xpc10nz) || (6'd37/*MS*/==-9'd245
              +xpc10nz) || (6'd37/*MS*/==-9'd244+xpc10nz) || (6'd37/*MS*/==-9'd242+xpc10nz) || (6'd37/*MS*/==-9'd241+xpc10nz) || (6'd37
              /*MS*/==-9'd239+xpc10nz) || (6'd37/*MS*/==-9'd238+xpc10nz) || (6'd37/*MS*/==-9'd236+xpc10nz) || (6'd37/*MS*/==-9'd171+xpc10nz
              ) || (6'd37/*MS*/==-8'd106+xpc10nz) || (6'd37/*MS*/==-8'd105+xpc10nz) || (6'd37/*MS*/==-8'd104+xpc10nz) || (6'd37/*MS*/==
              -8'd103+xpc10nz) || (6'd37/*MS*/==-8'd102+xpc10nz) || (6'd37/*MS*/==-8'd101+xpc10nz) || (6'd37/*MS*/==-8'd100+xpc10nz) || 
              (6'd37/*MS*/==-8'd99+xpc10nz) || (6'd37/*MS*/==-8'd98+xpc10nz) || (6'd37/*MS*/==-8'd97+xpc10nz) || (6'd37/*MS*/==-8'd96
              +xpc10nz) || (6'd37/*MS*/==-8'd95+xpc10nz) || (6'd37/*MS*/==-8'd94+xpc10nz) || (6'd37/*MS*/==-8'd93+xpc10nz) || (6'd37/*MS*/==
              -8'd92+xpc10nz) || (6'd37/*MS*/==-8'd91+xpc10nz) || (6'd37/*MS*/==-8'd90+xpc10nz) || (6'd37/*MS*/==-8'd89+xpc10nz) || (6'd37
              /*MS*/==-8'd88+xpc10nz) || (6'd37/*MS*/==-8'd87+xpc10nz) || (6'd37/*MS*/==-8'd86+xpc10nz) || (6'd37/*MS*/==-8'd85+xpc10nz
              ) || (6'd37/*MS*/==-8'd84+xpc10nz) || (6'd37/*MS*/==-8'd83+xpc10nz) || (6'd37/*MS*/==-8'd82+xpc10nz) || (6'd37/*MS*/==-8'd65
              +xpc10nz) || (6'd37/*MS*/==-8'd64+xpc10nz) || (6'd37/*MS*/==-7'd59+xpc10nz) || (6'd37/*MS*/==-7'd50+xpc10nz) || (6'd37/*MS*/==
              -7'd37+xpc10nz) || (6'd37/*MS*/==-6'd20+xpc10nz) || (6'd37/*MS*/==-6'd19+xpc10nz) || (6'd37/*MS*/==-6'd18+xpc10nz) || (6'd37
              /*MS*/==-6'd17+xpc10nz) || (6'd37/*MS*/==-6'd16+xpc10nz) || (6'd37/*MS*/==-5'd15+xpc10nz) || (6'd37/*MS*/==-5'd14+xpc10nz
              ) || (6'd37/*MS*/==-5'd13+xpc10nz) || (6'd37/*MS*/==-5'd12+xpc10nz) || (6'd37/*MS*/==-5'd11+xpc10nz) || (6'd37/*MS*/==-5'd10
              +xpc10nz) || (6'd37/*MS*/==-5'd9+xpc10nz) || (6'd37/*MS*/==-5'd8+xpc10nz) || (6'd37/*MS*/==-4'd7+xpc10nz) || (6'd37/*MS*/==
              -4'd6+xpc10nz) || (6'd37/*MS*/==-4'd5+xpc10nz) || (6'd37/*MS*/==-4'd4+xpc10nz) || (6'd37/*MS*/==-3'd3+xpc10nz) || (6'd37
              /*MS*/==-3'd2+xpc10nz) || (6'd37/*MS*/==-2'd1+xpc10nz) || (xpc10nz==6'd37/*US*/)) && !xpc10_clear && !xpc10_stall;

               xpc10_trk36 <= ((6'd36/*MS*/==-11'd609+xpc10nz) || (6'd36/*MS*/==-11'd599+xpc10nz) || (6'd36/*MS*/==-11'd588+xpc10nz) || 
              (6'd36/*MS*/==-11'd576+xpc10nz) || (6'd36/*MS*/==-11'd571+xpc10nz) || (6'd36/*MS*/==-11'd565+xpc10nz) || (6'd36/*MS*/==
              -11'd558+xpc10nz) || (6'd36/*MS*/==-11'd550+xpc10nz) || (6'd36/*MS*/==-11'd549+xpc10nz) || (6'd36/*MS*/==-11'd547+xpc10nz
              ) || (6'd36/*MS*/==-11'd544+xpc10nz) || (6'd36/*MS*/==-11'd540+xpc10nz) || (6'd36/*MS*/==-11'd539+xpc10nz) || (6'd36/*MS*/==
              -11'd537+xpc10nz) || (6'd36/*MS*/==-11'd534+xpc10nz) || (6'd36/*MS*/==-11'd532+xpc10nz) || (6'd36/*MS*/==-11'd528+xpc10nz
              ) || (6'd36/*MS*/==-10'd503+xpc10nz) || (6'd36/*MS*/==-10'd502+xpc10nz) || (6'd36/*MS*/==-10'd472+xpc10nz) || (6'd36/*MS*/==
              -10'd407+xpc10nz) || (6'd36/*MS*/==-10'd342+xpc10nz) || (6'd36/*MS*/==-10'd341+xpc10nz) || (6'd36/*MS*/==-10'd340+xpc10nz
              ) || (6'd36/*MS*/==-10'd338+xpc10nz) || (6'd36/*MS*/==-10'd335+xpc10nz) || (6'd36/*MS*/==-10'd334+xpc10nz) || (6'd36/*MS*/==
              -10'd330+xpc10nz) || (6'd36/*MS*/==-10'd329+xpc10nz) || (6'd36/*MS*/==-10'd327+xpc10nz) || (6'd36/*MS*/==-10'd324+xpc10nz
              ) || (6'd36/*MS*/==-10'd323+xpc10nz) || (6'd36/*MS*/==-10'd322+xpc10nz) || (6'd36/*MS*/==-10'd321+xpc10nz) || (6'd36/*MS*/==
              -10'd320+xpc10nz) || (6'd36/*MS*/==-10'd319+xpc10nz) || (6'd36/*MS*/==-10'd318+xpc10nz) || (6'd36/*MS*/==-10'd314+xpc10nz
              ) || (6'd36/*MS*/==-10'd289+xpc10nz) || (6'd36/*MS*/==-10'd287+xpc10nz) || (6'd36/*MS*/==-10'd285+xpc10nz) || (6'd36/*MS*/==
              -10'd284+xpc10nz) || (6'd36/*MS*/==-10'd259+xpc10nz) || (6'd36/*MS*/==-10'd258+xpc10nz) || (6'd36/*MS*/==-10'd257+xpc10nz
              ) || (6'd36/*MS*/==-9'd255+xpc10nz) || (6'd36/*MS*/==-9'd254+xpc10nz) || (6'd36/*MS*/==-9'd253+xpc10nz) || (6'd36/*MS*/==
              -9'd252+xpc10nz) || (6'd36/*MS*/==-9'd251+xpc10nz) || (6'd36/*MS*/==-9'd250+xpc10nz) || (6'd36/*MS*/==-9'd249+xpc10nz) || 
              (6'd36/*MS*/==-9'd248+xpc10nz) || (6'd36/*MS*/==-9'd247+xpc10nz) || (6'd36/*MS*/==-9'd246+xpc10nz) || (6'd36/*MS*/==-9'd245
              +xpc10nz) || (6'd36/*MS*/==-9'd244+xpc10nz) || (6'd36/*MS*/==-9'd242+xpc10nz) || (6'd36/*MS*/==-9'd241+xpc10nz) || (6'd36
              /*MS*/==-9'd239+xpc10nz) || (6'd36/*MS*/==-9'd238+xpc10nz) || (6'd36/*MS*/==-9'd236+xpc10nz) || (6'd36/*MS*/==-9'd171+xpc10nz
              ) || (6'd36/*MS*/==-8'd106+xpc10nz) || (6'd36/*MS*/==-8'd105+xpc10nz) || (6'd36/*MS*/==-8'd104+xpc10nz) || (6'd36/*MS*/==
              -8'd103+xpc10nz) || (6'd36/*MS*/==-8'd102+xpc10nz) || (6'd36/*MS*/==-8'd101+xpc10nz) || (6'd36/*MS*/==-8'd100+xpc10nz) || 
              (6'd36/*MS*/==-8'd99+xpc10nz) || (6'd36/*MS*/==-8'd98+xpc10nz) || (6'd36/*MS*/==-8'd97+xpc10nz) || (6'd36/*MS*/==-8'd96
              +xpc10nz) || (6'd36/*MS*/==-8'd95+xpc10nz) || (6'd36/*MS*/==-8'd94+xpc10nz) || (6'd36/*MS*/==-8'd93+xpc10nz) || (6'd36/*MS*/==
              -8'd92+xpc10nz) || (6'd36/*MS*/==-8'd91+xpc10nz) || (6'd36/*MS*/==-8'd90+xpc10nz) || (6'd36/*MS*/==-8'd89+xpc10nz) || (6'd36
              /*MS*/==-8'd88+xpc10nz) || (6'd36/*MS*/==-8'd87+xpc10nz) || (6'd36/*MS*/==-8'd86+xpc10nz) || (6'd36/*MS*/==-8'd85+xpc10nz
              ) || (6'd36/*MS*/==-8'd84+xpc10nz) || (6'd36/*MS*/==-8'd83+xpc10nz) || (6'd36/*MS*/==-8'd82+xpc10nz) || (6'd36/*MS*/==-8'd65
              +xpc10nz) || (6'd36/*MS*/==-8'd64+xpc10nz) || (6'd36/*MS*/==-7'd59+xpc10nz) || (6'd36/*MS*/==-7'd50+xpc10nz) || (6'd36/*MS*/==
              -7'd37+xpc10nz) || (6'd36/*MS*/==-6'd20+xpc10nz) || (6'd36/*MS*/==-6'd19+xpc10nz) || (6'd36/*MS*/==-6'd18+xpc10nz) || (6'd36
              /*MS*/==-6'd17+xpc10nz) || (6'd36/*MS*/==-6'd16+xpc10nz) || (6'd36/*MS*/==-5'd15+xpc10nz) || (6'd36/*MS*/==-5'd14+xpc10nz
              ) || (6'd36/*MS*/==-5'd13+xpc10nz) || (6'd36/*MS*/==-5'd12+xpc10nz) || (6'd36/*MS*/==-5'd11+xpc10nz) || (6'd36/*MS*/==-5'd10
              +xpc10nz) || (6'd36/*MS*/==-5'd9+xpc10nz) || (6'd36/*MS*/==-5'd8+xpc10nz) || (6'd36/*MS*/==-4'd7+xpc10nz) || (6'd36/*MS*/==
              -4'd6+xpc10nz) || (6'd36/*MS*/==-4'd5+xpc10nz) || (6'd36/*MS*/==-4'd4+xpc10nz) || (6'd36/*MS*/==-3'd3+xpc10nz) || (6'd36
              /*MS*/==-3'd2+xpc10nz) || (6'd36/*MS*/==-2'd1+xpc10nz) || (xpc10nz==6'd36/*US*/)) && !xpc10_clear && !xpc10_stall;

               xpc10_trk35 <= ((6'd35/*MS*/==-11'd609+xpc10nz) || (6'd35/*MS*/==-11'd599+xpc10nz) || (6'd35/*MS*/==-11'd588+xpc10nz) || 
              (6'd35/*MS*/==-11'd576+xpc10nz) || (6'd35/*MS*/==-11'd571+xpc10nz) || (6'd35/*MS*/==-11'd565+xpc10nz) || (6'd35/*MS*/==
              -11'd558+xpc10nz) || (6'd35/*MS*/==-11'd550+xpc10nz) || (6'd35/*MS*/==-11'd549+xpc10nz) || (6'd35/*MS*/==-11'd547+xpc10nz
              ) || (6'd35/*MS*/==-11'd544+xpc10nz) || (6'd35/*MS*/==-11'd540+xpc10nz) || (6'd35/*MS*/==-11'd539+xpc10nz) || (6'd35/*MS*/==
              -11'd537+xpc10nz) || (6'd35/*MS*/==-11'd534+xpc10nz) || (6'd35/*MS*/==-11'd532+xpc10nz) || (6'd35/*MS*/==-11'd528+xpc10nz
              ) || (6'd35/*MS*/==-10'd503+xpc10nz) || (6'd35/*MS*/==-10'd502+xpc10nz) || (6'd35/*MS*/==-10'd472+xpc10nz) || (6'd35/*MS*/==
              -10'd407+xpc10nz) || (6'd35/*MS*/==-10'd342+xpc10nz) || (6'd35/*MS*/==-10'd341+xpc10nz) || (6'd35/*MS*/==-10'd340+xpc10nz
              ) || (6'd35/*MS*/==-10'd338+xpc10nz) || (6'd35/*MS*/==-10'd335+xpc10nz) || (6'd35/*MS*/==-10'd334+xpc10nz) || (6'd35/*MS*/==
              -10'd330+xpc10nz) || (6'd35/*MS*/==-10'd329+xpc10nz) || (6'd35/*MS*/==-10'd327+xpc10nz) || (6'd35/*MS*/==-10'd324+xpc10nz
              ) || (6'd35/*MS*/==-10'd323+xpc10nz) || (6'd35/*MS*/==-10'd322+xpc10nz) || (6'd35/*MS*/==-10'd321+xpc10nz) || (6'd35/*MS*/==
              -10'd320+xpc10nz) || (6'd35/*MS*/==-10'd319+xpc10nz) || (6'd35/*MS*/==-10'd318+xpc10nz) || (6'd35/*MS*/==-10'd314+xpc10nz
              ) || (6'd35/*MS*/==-10'd289+xpc10nz) || (6'd35/*MS*/==-10'd287+xpc10nz) || (6'd35/*MS*/==-10'd285+xpc10nz) || (6'd35/*MS*/==
              -10'd284+xpc10nz) || (6'd35/*MS*/==-10'd259+xpc10nz) || (6'd35/*MS*/==-10'd258+xpc10nz) || (6'd35/*MS*/==-10'd257+xpc10nz
              ) || (6'd35/*MS*/==-9'd255+xpc10nz) || (6'd35/*MS*/==-9'd254+xpc10nz) || (6'd35/*MS*/==-9'd253+xpc10nz) || (6'd35/*MS*/==
              -9'd252+xpc10nz) || (6'd35/*MS*/==-9'd251+xpc10nz) || (6'd35/*MS*/==-9'd250+xpc10nz) || (6'd35/*MS*/==-9'd249+xpc10nz) || 
              (6'd35/*MS*/==-9'd248+xpc10nz) || (6'd35/*MS*/==-9'd247+xpc10nz) || (6'd35/*MS*/==-9'd246+xpc10nz) || (6'd35/*MS*/==-9'd245
              +xpc10nz) || (6'd35/*MS*/==-9'd244+xpc10nz) || (6'd35/*MS*/==-9'd242+xpc10nz) || (6'd35/*MS*/==-9'd241+xpc10nz) || (6'd35
              /*MS*/==-9'd239+xpc10nz) || (6'd35/*MS*/==-9'd238+xpc10nz) || (6'd35/*MS*/==-9'd236+xpc10nz) || (6'd35/*MS*/==-9'd171+xpc10nz
              ) || (6'd35/*MS*/==-8'd106+xpc10nz) || (6'd35/*MS*/==-8'd105+xpc10nz) || (6'd35/*MS*/==-8'd104+xpc10nz) || (6'd35/*MS*/==
              -8'd103+xpc10nz) || (6'd35/*MS*/==-8'd102+xpc10nz) || (6'd35/*MS*/==-8'd101+xpc10nz) || (6'd35/*MS*/==-8'd100+xpc10nz) || 
              (6'd35/*MS*/==-8'd99+xpc10nz) || (6'd35/*MS*/==-8'd98+xpc10nz) || (6'd35/*MS*/==-8'd97+xpc10nz) || (6'd35/*MS*/==-8'd96
              +xpc10nz) || (6'd35/*MS*/==-8'd95+xpc10nz) || (6'd35/*MS*/==-8'd94+xpc10nz) || (6'd35/*MS*/==-8'd93+xpc10nz) || (6'd35/*MS*/==
              -8'd92+xpc10nz) || (6'd35/*MS*/==-8'd91+xpc10nz) || (6'd35/*MS*/==-8'd90+xpc10nz) || (6'd35/*MS*/==-8'd89+xpc10nz) || (6'd35
              /*MS*/==-8'd88+xpc10nz) || (6'd35/*MS*/==-8'd87+xpc10nz) || (6'd35/*MS*/==-8'd86+xpc10nz) || (6'd35/*MS*/==-8'd85+xpc10nz
              ) || (6'd35/*MS*/==-8'd84+xpc10nz) || (6'd35/*MS*/==-8'd83+xpc10nz) || (6'd35/*MS*/==-8'd82+xpc10nz) || (6'd35/*MS*/==-8'd65
              +xpc10nz) || (6'd35/*MS*/==-8'd64+xpc10nz) || (6'd35/*MS*/==-7'd59+xpc10nz) || (6'd35/*MS*/==-7'd50+xpc10nz) || (6'd35/*MS*/==
              -7'd37+xpc10nz) || (6'd35/*MS*/==-6'd20+xpc10nz) || (6'd35/*MS*/==-6'd19+xpc10nz) || (6'd35/*MS*/==-6'd18+xpc10nz) || (6'd35
              /*MS*/==-6'd17+xpc10nz) || (6'd35/*MS*/==-6'd16+xpc10nz) || (6'd35/*MS*/==-5'd15+xpc10nz) || (6'd35/*MS*/==-5'd14+xpc10nz
              ) || (6'd35/*MS*/==-5'd13+xpc10nz) || (6'd35/*MS*/==-5'd12+xpc10nz) || (6'd35/*MS*/==-5'd11+xpc10nz) || (6'd35/*MS*/==-5'd10
              +xpc10nz) || (6'd35/*MS*/==-5'd9+xpc10nz) || (6'd35/*MS*/==-5'd8+xpc10nz) || (6'd35/*MS*/==-4'd7+xpc10nz) || (6'd35/*MS*/==
              -4'd6+xpc10nz) || (6'd35/*MS*/==-4'd5+xpc10nz) || (6'd35/*MS*/==-4'd4+xpc10nz) || (6'd35/*MS*/==-3'd3+xpc10nz) || (6'd35
              /*MS*/==-3'd2+xpc10nz) || (6'd35/*MS*/==-2'd1+xpc10nz) || (xpc10nz==6'd35/*US*/)) && !xpc10_clear && !xpc10_stall;

               xpc10_trk34 <= ((6'd34/*MS*/==-11'd609+xpc10nz) || (6'd34/*MS*/==-11'd599+xpc10nz) || (6'd34/*MS*/==-11'd588+xpc10nz) || 
              (6'd34/*MS*/==-11'd576+xpc10nz) || (6'd34/*MS*/==-11'd571+xpc10nz) || (6'd34/*MS*/==-11'd565+xpc10nz) || (6'd34/*MS*/==
              -11'd558+xpc10nz) || (6'd34/*MS*/==-11'd550+xpc10nz) || (6'd34/*MS*/==-11'd549+xpc10nz) || (6'd34/*MS*/==-11'd547+xpc10nz
              ) || (6'd34/*MS*/==-11'd544+xpc10nz) || (6'd34/*MS*/==-11'd540+xpc10nz) || (6'd34/*MS*/==-11'd539+xpc10nz) || (6'd34/*MS*/==
              -11'd537+xpc10nz) || (6'd34/*MS*/==-11'd534+xpc10nz) || (6'd34/*MS*/==-11'd532+xpc10nz) || (6'd34/*MS*/==-11'd528+xpc10nz
              ) || (6'd34/*MS*/==-10'd503+xpc10nz) || (6'd34/*MS*/==-10'd502+xpc10nz) || (6'd34/*MS*/==-10'd472+xpc10nz) || (6'd34/*MS*/==
              -10'd407+xpc10nz) || (6'd34/*MS*/==-10'd342+xpc10nz) || (6'd34/*MS*/==-10'd341+xpc10nz) || (6'd34/*MS*/==-10'd340+xpc10nz
              ) || (6'd34/*MS*/==-10'd338+xpc10nz) || (6'd34/*MS*/==-10'd335+xpc10nz) || (6'd34/*MS*/==-10'd334+xpc10nz) || (6'd34/*MS*/==
              -10'd330+xpc10nz) || (6'd34/*MS*/==-10'd329+xpc10nz) || (6'd34/*MS*/==-10'd327+xpc10nz) || (6'd34/*MS*/==-10'd324+xpc10nz
              ) || (6'd34/*MS*/==-10'd323+xpc10nz) || (6'd34/*MS*/==-10'd322+xpc10nz) || (6'd34/*MS*/==-10'd321+xpc10nz) || (6'd34/*MS*/==
              -10'd320+xpc10nz) || (6'd34/*MS*/==-10'd319+xpc10nz) || (6'd34/*MS*/==-10'd318+xpc10nz) || (6'd34/*MS*/==-10'd314+xpc10nz
              ) || (6'd34/*MS*/==-10'd289+xpc10nz) || (6'd34/*MS*/==-10'd287+xpc10nz) || (6'd34/*MS*/==-10'd285+xpc10nz) || (6'd34/*MS*/==
              -10'd284+xpc10nz) || (6'd34/*MS*/==-10'd259+xpc10nz) || (6'd34/*MS*/==-10'd258+xpc10nz) || (6'd34/*MS*/==-10'd257+xpc10nz
              ) || (6'd34/*MS*/==-9'd255+xpc10nz) || (6'd34/*MS*/==-9'd254+xpc10nz) || (6'd34/*MS*/==-9'd253+xpc10nz) || (6'd34/*MS*/==
              -9'd252+xpc10nz) || (6'd34/*MS*/==-9'd251+xpc10nz) || (6'd34/*MS*/==-9'd250+xpc10nz) || (6'd34/*MS*/==-9'd249+xpc10nz) || 
              (6'd34/*MS*/==-9'd248+xpc10nz) || (6'd34/*MS*/==-9'd247+xpc10nz) || (6'd34/*MS*/==-9'd246+xpc10nz) || (6'd34/*MS*/==-9'd245
              +xpc10nz) || (6'd34/*MS*/==-9'd244+xpc10nz) || (6'd34/*MS*/==-9'd242+xpc10nz) || (6'd34/*MS*/==-9'd241+xpc10nz) || (6'd34
              /*MS*/==-9'd239+xpc10nz) || (6'd34/*MS*/==-9'd238+xpc10nz) || (6'd34/*MS*/==-9'd236+xpc10nz) || (6'd34/*MS*/==-9'd171+xpc10nz
              ) || (6'd34/*MS*/==-8'd106+xpc10nz) || (6'd34/*MS*/==-8'd105+xpc10nz) || (6'd34/*MS*/==-8'd104+xpc10nz) || (6'd34/*MS*/==
              -8'd103+xpc10nz) || (6'd34/*MS*/==-8'd102+xpc10nz) || (6'd34/*MS*/==-8'd101+xpc10nz) || (6'd34/*MS*/==-8'd100+xpc10nz) || 
              (6'd34/*MS*/==-8'd99+xpc10nz) || (6'd34/*MS*/==-8'd98+xpc10nz) || (6'd34/*MS*/==-8'd97+xpc10nz) || (6'd34/*MS*/==-8'd96
              +xpc10nz) || (6'd34/*MS*/==-8'd95+xpc10nz) || (6'd34/*MS*/==-8'd94+xpc10nz) || (6'd34/*MS*/==-8'd93+xpc10nz) || (6'd34/*MS*/==
              -8'd92+xpc10nz) || (6'd34/*MS*/==-8'd91+xpc10nz) || (6'd34/*MS*/==-8'd90+xpc10nz) || (6'd34/*MS*/==-8'd89+xpc10nz) || (6'd34
              /*MS*/==-8'd88+xpc10nz) || (6'd34/*MS*/==-8'd87+xpc10nz) || (6'd34/*MS*/==-8'd86+xpc10nz) || (6'd34/*MS*/==-8'd85+xpc10nz
              ) || (6'd34/*MS*/==-8'd84+xpc10nz) || (6'd34/*MS*/==-8'd83+xpc10nz) || (6'd34/*MS*/==-8'd82+xpc10nz) || (6'd34/*MS*/==-8'd65
              +xpc10nz) || (6'd34/*MS*/==-8'd64+xpc10nz) || (6'd34/*MS*/==-7'd59+xpc10nz) || (6'd34/*MS*/==-7'd50+xpc10nz) || (6'd34/*MS*/==
              -7'd37+xpc10nz) || (6'd34/*MS*/==-6'd20+xpc10nz) || (6'd34/*MS*/==-6'd19+xpc10nz) || (6'd34/*MS*/==-6'd18+xpc10nz) || (6'd34
              /*MS*/==-6'd17+xpc10nz) || (6'd34/*MS*/==-6'd16+xpc10nz) || (6'd34/*MS*/==-5'd15+xpc10nz) || (6'd34/*MS*/==-5'd14+xpc10nz
              ) || (6'd34/*MS*/==-5'd13+xpc10nz) || (6'd34/*MS*/==-5'd12+xpc10nz) || (6'd34/*MS*/==-5'd11+xpc10nz) || (6'd34/*MS*/==-5'd10
              +xpc10nz) || (6'd34/*MS*/==-5'd9+xpc10nz) || (6'd34/*MS*/==-5'd8+xpc10nz) || (6'd34/*MS*/==-4'd7+xpc10nz) || (6'd34/*MS*/==
              -4'd6+xpc10nz) || (6'd34/*MS*/==-4'd5+xpc10nz) || (6'd34/*MS*/==-4'd4+xpc10nz) || (6'd34/*MS*/==-3'd3+xpc10nz) || (6'd34
              /*MS*/==-3'd2+xpc10nz) || (6'd34/*MS*/==-2'd1+xpc10nz) || (xpc10nz==6'd34/*US*/)) && !xpc10_clear && !xpc10_stall;

               xpc10_trk33 <= ((6'd33/*MS*/==-11'd609+xpc10nz) || (6'd33/*MS*/==-11'd599+xpc10nz) || (6'd33/*MS*/==-11'd588+xpc10nz) || 
              (6'd33/*MS*/==-11'd576+xpc10nz) || (6'd33/*MS*/==-11'd571+xpc10nz) || (6'd33/*MS*/==-11'd565+xpc10nz) || (6'd33/*MS*/==
              -11'd558+xpc10nz) || (6'd33/*MS*/==-11'd550+xpc10nz) || (6'd33/*MS*/==-11'd549+xpc10nz) || (6'd33/*MS*/==-11'd547+xpc10nz
              ) || (6'd33/*MS*/==-11'd544+xpc10nz) || (6'd33/*MS*/==-11'd540+xpc10nz) || (6'd33/*MS*/==-11'd539+xpc10nz) || (6'd33/*MS*/==
              -11'd537+xpc10nz) || (6'd33/*MS*/==-11'd534+xpc10nz) || (6'd33/*MS*/==-11'd532+xpc10nz) || (6'd33/*MS*/==-11'd528+xpc10nz
              ) || (6'd33/*MS*/==-10'd503+xpc10nz) || (6'd33/*MS*/==-10'd502+xpc10nz) || (6'd33/*MS*/==-10'd472+xpc10nz) || (6'd33/*MS*/==
              -10'd407+xpc10nz) || (6'd33/*MS*/==-10'd342+xpc10nz) || (6'd33/*MS*/==-10'd341+xpc10nz) || (6'd33/*MS*/==-10'd340+xpc10nz
              ) || (6'd33/*MS*/==-10'd338+xpc10nz) || (6'd33/*MS*/==-10'd335+xpc10nz) || (6'd33/*MS*/==-10'd334+xpc10nz) || (6'd33/*MS*/==
              -10'd330+xpc10nz) || (6'd33/*MS*/==-10'd329+xpc10nz) || (6'd33/*MS*/==-10'd327+xpc10nz) || (6'd33/*MS*/==-10'd324+xpc10nz
              ) || (6'd33/*MS*/==-10'd323+xpc10nz) || (6'd33/*MS*/==-10'd322+xpc10nz) || (6'd33/*MS*/==-10'd321+xpc10nz) || (6'd33/*MS*/==
              -10'd320+xpc10nz) || (6'd33/*MS*/==-10'd319+xpc10nz) || (6'd33/*MS*/==-10'd318+xpc10nz) || (6'd33/*MS*/==-10'd314+xpc10nz
              ) || (6'd33/*MS*/==-10'd289+xpc10nz) || (6'd33/*MS*/==-10'd287+xpc10nz) || (6'd33/*MS*/==-10'd285+xpc10nz) || (6'd33/*MS*/==
              -10'd284+xpc10nz) || (6'd33/*MS*/==-10'd259+xpc10nz) || (6'd33/*MS*/==-10'd258+xpc10nz) || (6'd33/*MS*/==-10'd257+xpc10nz
              ) || (6'd33/*MS*/==-9'd255+xpc10nz) || (6'd33/*MS*/==-9'd254+xpc10nz) || (6'd33/*MS*/==-9'd253+xpc10nz) || (6'd33/*MS*/==
              -9'd252+xpc10nz) || (6'd33/*MS*/==-9'd251+xpc10nz) || (6'd33/*MS*/==-9'd250+xpc10nz) || (6'd33/*MS*/==-9'd249+xpc10nz) || 
              (6'd33/*MS*/==-9'd248+xpc10nz) || (6'd33/*MS*/==-9'd247+xpc10nz) || (6'd33/*MS*/==-9'd246+xpc10nz) || (6'd33/*MS*/==-9'd245
              +xpc10nz) || (6'd33/*MS*/==-9'd244+xpc10nz) || (6'd33/*MS*/==-9'd242+xpc10nz) || (6'd33/*MS*/==-9'd241+xpc10nz) || (6'd33
              /*MS*/==-9'd239+xpc10nz) || (6'd33/*MS*/==-9'd238+xpc10nz) || (6'd33/*MS*/==-9'd236+xpc10nz) || (6'd33/*MS*/==-9'd171+xpc10nz
              ) || (6'd33/*MS*/==-8'd106+xpc10nz) || (6'd33/*MS*/==-8'd105+xpc10nz) || (6'd33/*MS*/==-8'd104+xpc10nz) || (6'd33/*MS*/==
              -8'd103+xpc10nz) || (6'd33/*MS*/==-8'd102+xpc10nz) || (6'd33/*MS*/==-8'd101+xpc10nz) || (6'd33/*MS*/==-8'd100+xpc10nz) || 
              (6'd33/*MS*/==-8'd99+xpc10nz) || (6'd33/*MS*/==-8'd98+xpc10nz) || (6'd33/*MS*/==-8'd97+xpc10nz) || (6'd33/*MS*/==-8'd96
              +xpc10nz) || (6'd33/*MS*/==-8'd95+xpc10nz) || (6'd33/*MS*/==-8'd94+xpc10nz) || (6'd33/*MS*/==-8'd93+xpc10nz) || (6'd33/*MS*/==
              -8'd92+xpc10nz) || (6'd33/*MS*/==-8'd91+xpc10nz) || (6'd33/*MS*/==-8'd90+xpc10nz) || (6'd33/*MS*/==-8'd89+xpc10nz) || (6'd33
              /*MS*/==-8'd88+xpc10nz) || (6'd33/*MS*/==-8'd87+xpc10nz) || (6'd33/*MS*/==-8'd86+xpc10nz) || (6'd33/*MS*/==-8'd85+xpc10nz
              ) || (6'd33/*MS*/==-8'd84+xpc10nz) || (6'd33/*MS*/==-8'd83+xpc10nz) || (6'd33/*MS*/==-8'd82+xpc10nz) || (6'd33/*MS*/==-8'd65
              +xpc10nz) || (6'd33/*MS*/==-8'd64+xpc10nz) || (6'd33/*MS*/==-7'd59+xpc10nz) || (6'd33/*MS*/==-7'd50+xpc10nz) || (6'd33/*MS*/==
              -7'd37+xpc10nz) || (6'd33/*MS*/==-6'd20+xpc10nz) || (6'd33/*MS*/==-6'd19+xpc10nz) || (6'd33/*MS*/==-6'd18+xpc10nz) || (6'd33
              /*MS*/==-6'd17+xpc10nz) || (6'd33/*MS*/==-6'd16+xpc10nz) || (6'd33/*MS*/==-5'd15+xpc10nz) || (6'd33/*MS*/==-5'd14+xpc10nz
              ) || (6'd33/*MS*/==-5'd13+xpc10nz) || (6'd33/*MS*/==-5'd12+xpc10nz) || (6'd33/*MS*/==-5'd11+xpc10nz) || (6'd33/*MS*/==-5'd10
              +xpc10nz) || (6'd33/*MS*/==-5'd9+xpc10nz) || (6'd33/*MS*/==-5'd8+xpc10nz) || (6'd33/*MS*/==-4'd7+xpc10nz) || (6'd33/*MS*/==
              -4'd6+xpc10nz) || (6'd33/*MS*/==-4'd5+xpc10nz) || (6'd33/*MS*/==-4'd4+xpc10nz) || (6'd33/*MS*/==-3'd3+xpc10nz) || (6'd33
              /*MS*/==-3'd2+xpc10nz) || (6'd33/*MS*/==-2'd1+xpc10nz) || (xpc10nz==6'd33/*US*/)) && !xpc10_clear && !xpc10_stall;

               xpc10_trk32 <= ((6'd32/*MS*/==-11'd609+xpc10nz) || (6'd32/*MS*/==-11'd599+xpc10nz) || (6'd32/*MS*/==-11'd588+xpc10nz) || 
              (6'd32/*MS*/==-11'd576+xpc10nz) || (6'd32/*MS*/==-11'd571+xpc10nz) || (6'd32/*MS*/==-11'd565+xpc10nz) || (6'd32/*MS*/==
              -11'd558+xpc10nz) || (6'd32/*MS*/==-11'd550+xpc10nz) || (6'd32/*MS*/==-11'd549+xpc10nz) || (6'd32/*MS*/==-11'd547+xpc10nz
              ) || (6'd32/*MS*/==-11'd544+xpc10nz) || (6'd32/*MS*/==-11'd540+xpc10nz) || (6'd32/*MS*/==-11'd539+xpc10nz) || (6'd32/*MS*/==
              -11'd537+xpc10nz) || (6'd32/*MS*/==-11'd534+xpc10nz) || (6'd32/*MS*/==-11'd532+xpc10nz) || (6'd32/*MS*/==-11'd528+xpc10nz
              ) || (6'd32/*MS*/==-10'd503+xpc10nz) || (6'd32/*MS*/==-10'd502+xpc10nz) || (6'd32/*MS*/==-10'd472+xpc10nz) || (6'd32/*MS*/==
              -10'd407+xpc10nz) || (6'd32/*MS*/==-10'd342+xpc10nz) || (6'd32/*MS*/==-10'd341+xpc10nz) || (6'd32/*MS*/==-10'd340+xpc10nz
              ) || (6'd32/*MS*/==-10'd338+xpc10nz) || (6'd32/*MS*/==-10'd335+xpc10nz) || (6'd32/*MS*/==-10'd334+xpc10nz) || (6'd32/*MS*/==
              -10'd330+xpc10nz) || (6'd32/*MS*/==-10'd329+xpc10nz) || (6'd32/*MS*/==-10'd327+xpc10nz) || (6'd32/*MS*/==-10'd324+xpc10nz
              ) || (6'd32/*MS*/==-10'd323+xpc10nz) || (6'd32/*MS*/==-10'd322+xpc10nz) || (6'd32/*MS*/==-10'd321+xpc10nz) || (6'd32/*MS*/==
              -10'd320+xpc10nz) || (6'd32/*MS*/==-10'd319+xpc10nz) || (6'd32/*MS*/==-10'd318+xpc10nz) || (6'd32/*MS*/==-10'd314+xpc10nz
              ) || (6'd32/*MS*/==-10'd289+xpc10nz) || (6'd32/*MS*/==-10'd287+xpc10nz) || (6'd32/*MS*/==-10'd285+xpc10nz) || (6'd32/*MS*/==
              -10'd284+xpc10nz) || (6'd32/*MS*/==-10'd259+xpc10nz) || (6'd32/*MS*/==-10'd258+xpc10nz) || (6'd32/*MS*/==-10'd257+xpc10nz
              ) || (6'd32/*MS*/==-9'd255+xpc10nz) || (6'd32/*MS*/==-9'd254+xpc10nz) || (6'd32/*MS*/==-9'd253+xpc10nz) || (6'd32/*MS*/==
              -9'd252+xpc10nz) || (6'd32/*MS*/==-9'd251+xpc10nz) || (6'd32/*MS*/==-9'd250+xpc10nz) || (6'd32/*MS*/==-9'd249+xpc10nz) || 
              (6'd32/*MS*/==-9'd248+xpc10nz) || (6'd32/*MS*/==-9'd247+xpc10nz) || (6'd32/*MS*/==-9'd246+xpc10nz) || (6'd32/*MS*/==-9'd245
              +xpc10nz) || (6'd32/*MS*/==-9'd244+xpc10nz) || (6'd32/*MS*/==-9'd242+xpc10nz) || (6'd32/*MS*/==-9'd241+xpc10nz) || (6'd32
              /*MS*/==-9'd239+xpc10nz) || (6'd32/*MS*/==-9'd238+xpc10nz) || (6'd32/*MS*/==-9'd236+xpc10nz) || (6'd32/*MS*/==-9'd171+xpc10nz
              ) || (6'd32/*MS*/==-8'd106+xpc10nz) || (6'd32/*MS*/==-8'd105+xpc10nz) || (6'd32/*MS*/==-8'd104+xpc10nz) || (6'd32/*MS*/==
              -8'd103+xpc10nz) || (6'd32/*MS*/==-8'd102+xpc10nz) || (6'd32/*MS*/==-8'd101+xpc10nz) || (6'd32/*MS*/==-8'd100+xpc10nz) || 
              (6'd32/*MS*/==-8'd99+xpc10nz) || (6'd32/*MS*/==-8'd98+xpc10nz) || (6'd32/*MS*/==-8'd97+xpc10nz) || (6'd32/*MS*/==-8'd96
              +xpc10nz) || (6'd32/*MS*/==-8'd95+xpc10nz) || (6'd32/*MS*/==-8'd94+xpc10nz) || (6'd32/*MS*/==-8'd93+xpc10nz) || (6'd32/*MS*/==
              -8'd92+xpc10nz) || (6'd32/*MS*/==-8'd91+xpc10nz) || (6'd32/*MS*/==-8'd90+xpc10nz) || (6'd32/*MS*/==-8'd89+xpc10nz) || (6'd32
              /*MS*/==-8'd88+xpc10nz) || (6'd32/*MS*/==-8'd87+xpc10nz) || (6'd32/*MS*/==-8'd86+xpc10nz) || (6'd32/*MS*/==-8'd85+xpc10nz
              ) || (6'd32/*MS*/==-8'd84+xpc10nz) || (6'd32/*MS*/==-8'd83+xpc10nz) || (6'd32/*MS*/==-8'd82+xpc10nz) || (6'd32/*MS*/==-8'd65
              +xpc10nz) || (6'd32/*MS*/==-8'd64+xpc10nz) || (6'd32/*MS*/==-7'd59+xpc10nz) || (6'd32/*MS*/==-7'd50+xpc10nz) || (6'd32/*MS*/==
              -7'd37+xpc10nz) || (6'd32/*MS*/==-6'd20+xpc10nz) || (6'd32/*MS*/==-6'd19+xpc10nz) || (6'd32/*MS*/==-6'd18+xpc10nz) || (6'd32
              /*MS*/==-6'd17+xpc10nz) || (6'd32/*MS*/==-6'd16+xpc10nz) || (6'd32/*MS*/==-5'd15+xpc10nz) || (6'd32/*MS*/==-5'd14+xpc10nz
              ) || (6'd32/*MS*/==-5'd13+xpc10nz) || (6'd32/*MS*/==-5'd12+xpc10nz) || (6'd32/*MS*/==-5'd11+xpc10nz) || (6'd32/*MS*/==-5'd10
              +xpc10nz) || (6'd32/*MS*/==-5'd9+xpc10nz) || (6'd32/*MS*/==-5'd8+xpc10nz) || (6'd32/*MS*/==-4'd7+xpc10nz) || (6'd32/*MS*/==
              -4'd6+xpc10nz) || (6'd32/*MS*/==-4'd5+xpc10nz) || (6'd32/*MS*/==-4'd4+xpc10nz) || (6'd32/*MS*/==-3'd3+xpc10nz) || (6'd32
              /*MS*/==-3'd2+xpc10nz) || (6'd32/*MS*/==-2'd1+xpc10nz) || (xpc10nz==6'd32/*US*/)) && !xpc10_clear && !xpc10_stall;

               xpc10_trk31 <= ((5'd31/*MS*/==-11'd609+xpc10nz) || (5'd31/*MS*/==-11'd599+xpc10nz) || (5'd31/*MS*/==-11'd588+xpc10nz) || 
              (5'd31/*MS*/==-11'd576+xpc10nz) || (5'd31/*MS*/==-11'd571+xpc10nz) || (5'd31/*MS*/==-11'd565+xpc10nz) || (5'd31/*MS*/==
              -11'd558+xpc10nz) || (5'd31/*MS*/==-11'd550+xpc10nz) || (5'd31/*MS*/==-11'd549+xpc10nz) || (5'd31/*MS*/==-11'd547+xpc10nz
              ) || (5'd31/*MS*/==-11'd544+xpc10nz) || (5'd31/*MS*/==-11'd540+xpc10nz) || (5'd31/*MS*/==-11'd539+xpc10nz) || (5'd31/*MS*/==
              -11'd537+xpc10nz) || (5'd31/*MS*/==-11'd534+xpc10nz) || (5'd31/*MS*/==-11'd532+xpc10nz) || (5'd31/*MS*/==-11'd528+xpc10nz
              ) || (5'd31/*MS*/==-10'd503+xpc10nz) || (5'd31/*MS*/==-10'd502+xpc10nz) || (5'd31/*MS*/==-10'd472+xpc10nz) || (5'd31/*MS*/==
              -10'd407+xpc10nz) || (5'd31/*MS*/==-10'd342+xpc10nz) || (5'd31/*MS*/==-10'd341+xpc10nz) || (5'd31/*MS*/==-10'd340+xpc10nz
              ) || (5'd31/*MS*/==-10'd338+xpc10nz) || (5'd31/*MS*/==-10'd335+xpc10nz) || (5'd31/*MS*/==-10'd334+xpc10nz) || (5'd31/*MS*/==
              -10'd330+xpc10nz) || (5'd31/*MS*/==-10'd329+xpc10nz) || (5'd31/*MS*/==-10'd327+xpc10nz) || (5'd31/*MS*/==-10'd324+xpc10nz
              ) || (5'd31/*MS*/==-10'd323+xpc10nz) || (5'd31/*MS*/==-10'd322+xpc10nz) || (5'd31/*MS*/==-10'd321+xpc10nz) || (5'd31/*MS*/==
              -10'd320+xpc10nz) || (5'd31/*MS*/==-10'd319+xpc10nz) || (5'd31/*MS*/==-10'd318+xpc10nz) || (5'd31/*MS*/==-10'd314+xpc10nz
              ) || (5'd31/*MS*/==-10'd289+xpc10nz) || (5'd31/*MS*/==-10'd287+xpc10nz) || (5'd31/*MS*/==-10'd285+xpc10nz) || (5'd31/*MS*/==
              -10'd284+xpc10nz) || (5'd31/*MS*/==-10'd259+xpc10nz) || (5'd31/*MS*/==-10'd258+xpc10nz) || (5'd31/*MS*/==-10'd257+xpc10nz
              ) || (5'd31/*MS*/==-9'd255+xpc10nz) || (5'd31/*MS*/==-9'd254+xpc10nz) || (5'd31/*MS*/==-9'd253+xpc10nz) || (5'd31/*MS*/==
              -9'd252+xpc10nz) || (5'd31/*MS*/==-9'd251+xpc10nz) || (5'd31/*MS*/==-9'd250+xpc10nz) || (5'd31/*MS*/==-9'd249+xpc10nz) || 
              (5'd31/*MS*/==-9'd248+xpc10nz) || (5'd31/*MS*/==-9'd247+xpc10nz) || (5'd31/*MS*/==-9'd246+xpc10nz) || (5'd31/*MS*/==-9'd245
              +xpc10nz) || (5'd31/*MS*/==-9'd244+xpc10nz) || (5'd31/*MS*/==-9'd242+xpc10nz) || (5'd31/*MS*/==-9'd241+xpc10nz) || (5'd31
              /*MS*/==-9'd239+xpc10nz) || (5'd31/*MS*/==-9'd238+xpc10nz) || (5'd31/*MS*/==-9'd236+xpc10nz) || (5'd31/*MS*/==-9'd171+xpc10nz
              ) || (5'd31/*MS*/==-8'd106+xpc10nz) || (5'd31/*MS*/==-8'd105+xpc10nz) || (5'd31/*MS*/==-8'd104+xpc10nz) || (5'd31/*MS*/==
              -8'd103+xpc10nz) || (5'd31/*MS*/==-8'd102+xpc10nz) || (5'd31/*MS*/==-8'd101+xpc10nz) || (5'd31/*MS*/==-8'd100+xpc10nz) || 
              (5'd31/*MS*/==-8'd99+xpc10nz) || (5'd31/*MS*/==-8'd98+xpc10nz) || (5'd31/*MS*/==-8'd97+xpc10nz) || (5'd31/*MS*/==-8'd96
              +xpc10nz) || (5'd31/*MS*/==-8'd95+xpc10nz) || (5'd31/*MS*/==-8'd94+xpc10nz) || (5'd31/*MS*/==-8'd93+xpc10nz) || (5'd31/*MS*/==
              -8'd92+xpc10nz) || (5'd31/*MS*/==-8'd91+xpc10nz) || (5'd31/*MS*/==-8'd90+xpc10nz) || (5'd31/*MS*/==-8'd89+xpc10nz) || (5'd31
              /*MS*/==-8'd88+xpc10nz) || (5'd31/*MS*/==-8'd87+xpc10nz) || (5'd31/*MS*/==-8'd86+xpc10nz) || (5'd31/*MS*/==-8'd85+xpc10nz
              ) || (5'd31/*MS*/==-8'd84+xpc10nz) || (5'd31/*MS*/==-8'd83+xpc10nz) || (5'd31/*MS*/==-8'd82+xpc10nz) || (5'd31/*MS*/==-8'd65
              +xpc10nz) || (5'd31/*MS*/==-8'd64+xpc10nz) || (5'd31/*MS*/==-7'd59+xpc10nz) || (5'd31/*MS*/==-7'd50+xpc10nz) || (5'd31/*MS*/==
              -7'd37+xpc10nz) || (5'd31/*MS*/==-6'd20+xpc10nz) || (5'd31/*MS*/==-6'd19+xpc10nz) || (5'd31/*MS*/==-6'd18+xpc10nz) || (5'd31
              /*MS*/==-6'd17+xpc10nz) || (5'd31/*MS*/==-6'd16+xpc10nz) || (5'd31/*MS*/==-5'd15+xpc10nz) || (5'd31/*MS*/==-5'd14+xpc10nz
              ) || (5'd31/*MS*/==-5'd13+xpc10nz) || (5'd31/*MS*/==-5'd12+xpc10nz) || (5'd31/*MS*/==-5'd11+xpc10nz) || (5'd31/*MS*/==-5'd10
              +xpc10nz) || (5'd31/*MS*/==-5'd9+xpc10nz) || (5'd31/*MS*/==-5'd8+xpc10nz) || (5'd31/*MS*/==-4'd7+xpc10nz) || (5'd31/*MS*/==
              -4'd6+xpc10nz) || (5'd31/*MS*/==-4'd5+xpc10nz) || (5'd31/*MS*/==-4'd4+xpc10nz) || (5'd31/*MS*/==-3'd3+xpc10nz) || (5'd31
              /*MS*/==-3'd2+xpc10nz) || (5'd31/*MS*/==-2'd1+xpc10nz) || (xpc10nz==5'd31/*US*/)) && !xpc10_clear && !xpc10_stall;

               xpc10_trk30 <= ((5'd30/*MS*/==-11'd609+xpc10nz) || (5'd30/*MS*/==-11'd599+xpc10nz) || (5'd30/*MS*/==-11'd588+xpc10nz) || 
              (5'd30/*MS*/==-11'd576+xpc10nz) || (5'd30/*MS*/==-11'd571+xpc10nz) || (5'd30/*MS*/==-11'd565+xpc10nz) || (5'd30/*MS*/==
              -11'd558+xpc10nz) || (5'd30/*MS*/==-11'd550+xpc10nz) || (5'd30/*MS*/==-11'd549+xpc10nz) || (5'd30/*MS*/==-11'd547+xpc10nz
              ) || (5'd30/*MS*/==-11'd544+xpc10nz) || (5'd30/*MS*/==-11'd540+xpc10nz) || (5'd30/*MS*/==-11'd539+xpc10nz) || (5'd30/*MS*/==
              -11'd537+xpc10nz) || (5'd30/*MS*/==-11'd534+xpc10nz) || (5'd30/*MS*/==-11'd532+xpc10nz) || (5'd30/*MS*/==-11'd528+xpc10nz
              ) || (5'd30/*MS*/==-10'd503+xpc10nz) || (5'd30/*MS*/==-10'd502+xpc10nz) || (5'd30/*MS*/==-10'd472+xpc10nz) || (5'd30/*MS*/==
              -10'd407+xpc10nz) || (5'd30/*MS*/==-10'd342+xpc10nz) || (5'd30/*MS*/==-10'd341+xpc10nz) || (5'd30/*MS*/==-10'd340+xpc10nz
              ) || (5'd30/*MS*/==-10'd338+xpc10nz) || (5'd30/*MS*/==-10'd335+xpc10nz) || (5'd30/*MS*/==-10'd334+xpc10nz) || (5'd30/*MS*/==
              -10'd330+xpc10nz) || (5'd30/*MS*/==-10'd329+xpc10nz) || (5'd30/*MS*/==-10'd327+xpc10nz) || (5'd30/*MS*/==-10'd324+xpc10nz
              ) || (5'd30/*MS*/==-10'd323+xpc10nz) || (5'd30/*MS*/==-10'd322+xpc10nz) || (5'd30/*MS*/==-10'd321+xpc10nz) || (5'd30/*MS*/==
              -10'd320+xpc10nz) || (5'd30/*MS*/==-10'd319+xpc10nz) || (5'd30/*MS*/==-10'd318+xpc10nz) || (5'd30/*MS*/==-10'd314+xpc10nz
              ) || (5'd30/*MS*/==-10'd289+xpc10nz) || (5'd30/*MS*/==-10'd287+xpc10nz) || (5'd30/*MS*/==-10'd285+xpc10nz) || (5'd30/*MS*/==
              -10'd284+xpc10nz) || (5'd30/*MS*/==-10'd259+xpc10nz) || (5'd30/*MS*/==-10'd258+xpc10nz) || (5'd30/*MS*/==-10'd257+xpc10nz
              ) || (5'd30/*MS*/==-9'd255+xpc10nz) || (5'd30/*MS*/==-9'd254+xpc10nz) || (5'd30/*MS*/==-9'd253+xpc10nz) || (5'd30/*MS*/==
              -9'd252+xpc10nz) || (5'd30/*MS*/==-9'd251+xpc10nz) || (5'd30/*MS*/==-9'd250+xpc10nz) || (5'd30/*MS*/==-9'd249+xpc10nz) || 
              (5'd30/*MS*/==-9'd248+xpc10nz) || (5'd30/*MS*/==-9'd247+xpc10nz) || (5'd30/*MS*/==-9'd246+xpc10nz) || (5'd30/*MS*/==-9'd245
              +xpc10nz) || (5'd30/*MS*/==-9'd244+xpc10nz) || (5'd30/*MS*/==-9'd242+xpc10nz) || (5'd30/*MS*/==-9'd241+xpc10nz) || (5'd30
              /*MS*/==-9'd239+xpc10nz) || (5'd30/*MS*/==-9'd238+xpc10nz) || (5'd30/*MS*/==-9'd236+xpc10nz) || (5'd30/*MS*/==-9'd171+xpc10nz
              ) || (5'd30/*MS*/==-8'd106+xpc10nz) || (5'd30/*MS*/==-8'd105+xpc10nz) || (5'd30/*MS*/==-8'd104+xpc10nz) || (5'd30/*MS*/==
              -8'd103+xpc10nz) || (5'd30/*MS*/==-8'd102+xpc10nz) || (5'd30/*MS*/==-8'd101+xpc10nz) || (5'd30/*MS*/==-8'd100+xpc10nz) || 
              (5'd30/*MS*/==-8'd99+xpc10nz) || (5'd30/*MS*/==-8'd98+xpc10nz) || (5'd30/*MS*/==-8'd97+xpc10nz) || (5'd30/*MS*/==-8'd96
              +xpc10nz) || (5'd30/*MS*/==-8'd95+xpc10nz) || (5'd30/*MS*/==-8'd94+xpc10nz) || (5'd30/*MS*/==-8'd93+xpc10nz) || (5'd30/*MS*/==
              -8'd92+xpc10nz) || (5'd30/*MS*/==-8'd91+xpc10nz) || (5'd30/*MS*/==-8'd90+xpc10nz) || (5'd30/*MS*/==-8'd89+xpc10nz) || (5'd30
              /*MS*/==-8'd88+xpc10nz) || (5'd30/*MS*/==-8'd87+xpc10nz) || (5'd30/*MS*/==-8'd86+xpc10nz) || (5'd30/*MS*/==-8'd85+xpc10nz
              ) || (5'd30/*MS*/==-8'd84+xpc10nz) || (5'd30/*MS*/==-8'd83+xpc10nz) || (5'd30/*MS*/==-8'd82+xpc10nz) || (5'd30/*MS*/==-8'd65
              +xpc10nz) || (5'd30/*MS*/==-8'd64+xpc10nz) || (5'd30/*MS*/==-7'd59+xpc10nz) || (5'd30/*MS*/==-7'd50+xpc10nz) || (5'd30/*MS*/==
              -7'd37+xpc10nz) || (5'd30/*MS*/==-6'd20+xpc10nz) || (5'd30/*MS*/==-6'd19+xpc10nz) || (5'd30/*MS*/==-6'd18+xpc10nz) || (5'd30
              /*MS*/==-6'd17+xpc10nz) || (5'd30/*MS*/==-6'd16+xpc10nz) || (5'd30/*MS*/==-5'd15+xpc10nz) || (5'd30/*MS*/==-5'd14+xpc10nz
              ) || (5'd30/*MS*/==-5'd13+xpc10nz) || (5'd30/*MS*/==-5'd12+xpc10nz) || (5'd30/*MS*/==-5'd11+xpc10nz) || (5'd30/*MS*/==-5'd10
              +xpc10nz) || (5'd30/*MS*/==-5'd9+xpc10nz) || (5'd30/*MS*/==-5'd8+xpc10nz) || (5'd30/*MS*/==-4'd7+xpc10nz) || (5'd30/*MS*/==
              -4'd6+xpc10nz) || (5'd30/*MS*/==-4'd5+xpc10nz) || (5'd30/*MS*/==-4'd4+xpc10nz) || (5'd30/*MS*/==-3'd3+xpc10nz) || (5'd30
              /*MS*/==-3'd2+xpc10nz) || (5'd30/*MS*/==-2'd1+xpc10nz) || (xpc10nz==5'd30/*US*/)) && !xpc10_clear && !xpc10_stall;

               xpc10_trk29 <= ((5'd29/*MS*/==-11'd609+xpc10nz) || (5'd29/*MS*/==-11'd599+xpc10nz) || (5'd29/*MS*/==-11'd588+xpc10nz) || 
              (5'd29/*MS*/==-11'd576+xpc10nz) || (5'd29/*MS*/==-11'd571+xpc10nz) || (5'd29/*MS*/==-11'd565+xpc10nz) || (5'd29/*MS*/==
              -11'd558+xpc10nz) || (5'd29/*MS*/==-11'd550+xpc10nz) || (5'd29/*MS*/==-11'd549+xpc10nz) || (5'd29/*MS*/==-11'd547+xpc10nz
              ) || (5'd29/*MS*/==-11'd544+xpc10nz) || (5'd29/*MS*/==-11'd540+xpc10nz) || (5'd29/*MS*/==-11'd539+xpc10nz) || (5'd29/*MS*/==
              -11'd537+xpc10nz) || (5'd29/*MS*/==-11'd534+xpc10nz) || (5'd29/*MS*/==-11'd532+xpc10nz) || (5'd29/*MS*/==-11'd528+xpc10nz
              ) || (5'd29/*MS*/==-10'd503+xpc10nz) || (5'd29/*MS*/==-10'd502+xpc10nz) || (5'd29/*MS*/==-10'd472+xpc10nz) || (5'd29/*MS*/==
              -10'd407+xpc10nz) || (5'd29/*MS*/==-10'd342+xpc10nz) || (5'd29/*MS*/==-10'd341+xpc10nz) || (5'd29/*MS*/==-10'd340+xpc10nz
              ) || (5'd29/*MS*/==-10'd338+xpc10nz) || (5'd29/*MS*/==-10'd335+xpc10nz) || (5'd29/*MS*/==-10'd334+xpc10nz) || (5'd29/*MS*/==
              -10'd330+xpc10nz) || (5'd29/*MS*/==-10'd329+xpc10nz) || (5'd29/*MS*/==-10'd327+xpc10nz) || (5'd29/*MS*/==-10'd324+xpc10nz
              ) || (5'd29/*MS*/==-10'd323+xpc10nz) || (5'd29/*MS*/==-10'd322+xpc10nz) || (5'd29/*MS*/==-10'd321+xpc10nz) || (5'd29/*MS*/==
              -10'd320+xpc10nz) || (5'd29/*MS*/==-10'd319+xpc10nz) || (5'd29/*MS*/==-10'd318+xpc10nz) || (5'd29/*MS*/==-10'd314+xpc10nz
              ) || (5'd29/*MS*/==-10'd289+xpc10nz) || (5'd29/*MS*/==-10'd287+xpc10nz) || (5'd29/*MS*/==-10'd285+xpc10nz) || (5'd29/*MS*/==
              -10'd284+xpc10nz) || (5'd29/*MS*/==-10'd259+xpc10nz) || (5'd29/*MS*/==-10'd258+xpc10nz) || (5'd29/*MS*/==-10'd257+xpc10nz
              ) || (5'd29/*MS*/==-9'd255+xpc10nz) || (5'd29/*MS*/==-9'd254+xpc10nz) || (5'd29/*MS*/==-9'd253+xpc10nz) || (5'd29/*MS*/==
              -9'd252+xpc10nz) || (5'd29/*MS*/==-9'd251+xpc10nz) || (5'd29/*MS*/==-9'd250+xpc10nz) || (5'd29/*MS*/==-9'd249+xpc10nz) || 
              (5'd29/*MS*/==-9'd248+xpc10nz) || (5'd29/*MS*/==-9'd247+xpc10nz) || (5'd29/*MS*/==-9'd246+xpc10nz) || (5'd29/*MS*/==-9'd245
              +xpc10nz) || (5'd29/*MS*/==-9'd244+xpc10nz) || (5'd29/*MS*/==-9'd242+xpc10nz) || (5'd29/*MS*/==-9'd241+xpc10nz) || (5'd29
              /*MS*/==-9'd239+xpc10nz) || (5'd29/*MS*/==-9'd238+xpc10nz) || (5'd29/*MS*/==-9'd236+xpc10nz) || (5'd29/*MS*/==-9'd171+xpc10nz
              ) || (5'd29/*MS*/==-8'd106+xpc10nz) || (5'd29/*MS*/==-8'd105+xpc10nz) || (5'd29/*MS*/==-8'd104+xpc10nz) || (5'd29/*MS*/==
              -8'd103+xpc10nz) || (5'd29/*MS*/==-8'd102+xpc10nz) || (5'd29/*MS*/==-8'd101+xpc10nz) || (5'd29/*MS*/==-8'd100+xpc10nz) || 
              (5'd29/*MS*/==-8'd99+xpc10nz) || (5'd29/*MS*/==-8'd98+xpc10nz) || (5'd29/*MS*/==-8'd97+xpc10nz) || (5'd29/*MS*/==-8'd96
              +xpc10nz) || (5'd29/*MS*/==-8'd95+xpc10nz) || (5'd29/*MS*/==-8'd94+xpc10nz) || (5'd29/*MS*/==-8'd93+xpc10nz) || (5'd29/*MS*/==
              -8'd92+xpc10nz) || (5'd29/*MS*/==-8'd91+xpc10nz) || (5'd29/*MS*/==-8'd90+xpc10nz) || (5'd29/*MS*/==-8'd89+xpc10nz) || (5'd29
              /*MS*/==-8'd88+xpc10nz) || (5'd29/*MS*/==-8'd87+xpc10nz) || (5'd29/*MS*/==-8'd86+xpc10nz) || (5'd29/*MS*/==-8'd85+xpc10nz
              ) || (5'd29/*MS*/==-8'd84+xpc10nz) || (5'd29/*MS*/==-8'd83+xpc10nz) || (5'd29/*MS*/==-8'd82+xpc10nz) || (5'd29/*MS*/==-8'd65
              +xpc10nz) || (5'd29/*MS*/==-8'd64+xpc10nz) || (5'd29/*MS*/==-7'd59+xpc10nz) || (5'd29/*MS*/==-7'd50+xpc10nz) || (5'd29/*MS*/==
              -7'd37+xpc10nz) || (5'd29/*MS*/==-6'd20+xpc10nz) || (5'd29/*MS*/==-6'd19+xpc10nz) || (5'd29/*MS*/==-6'd18+xpc10nz) || (5'd29
              /*MS*/==-6'd17+xpc10nz) || (5'd29/*MS*/==-6'd16+xpc10nz) || (5'd29/*MS*/==-5'd15+xpc10nz) || (5'd29/*MS*/==-5'd14+xpc10nz
              ) || (5'd29/*MS*/==-5'd13+xpc10nz) || (5'd29/*MS*/==-5'd12+xpc10nz) || (5'd29/*MS*/==-5'd11+xpc10nz) || (5'd29/*MS*/==-5'd10
              +xpc10nz) || (5'd29/*MS*/==-5'd9+xpc10nz) || (5'd29/*MS*/==-5'd8+xpc10nz) || (5'd29/*MS*/==-4'd7+xpc10nz) || (5'd29/*MS*/==
              -4'd6+xpc10nz) || (5'd29/*MS*/==-4'd5+xpc10nz) || (5'd29/*MS*/==-4'd4+xpc10nz) || (5'd29/*MS*/==-3'd3+xpc10nz) || (5'd29
              /*MS*/==-3'd2+xpc10nz) || (5'd29/*MS*/==-2'd1+xpc10nz) || (xpc10nz==5'd29/*US*/)) && !xpc10_clear && !xpc10_stall;

               xpc10_trk28 <= ((5'd28/*MS*/==-11'd609+xpc10nz) || (5'd28/*MS*/==-11'd599+xpc10nz) || (5'd28/*MS*/==-11'd588+xpc10nz) || 
              (5'd28/*MS*/==-11'd576+xpc10nz) || (5'd28/*MS*/==-11'd571+xpc10nz) || (5'd28/*MS*/==-11'd565+xpc10nz) || (5'd28/*MS*/==
              -11'd558+xpc10nz) || (5'd28/*MS*/==-11'd550+xpc10nz) || (5'd28/*MS*/==-11'd549+xpc10nz) || (5'd28/*MS*/==-11'd547+xpc10nz
              ) || (5'd28/*MS*/==-11'd544+xpc10nz) || (5'd28/*MS*/==-11'd540+xpc10nz) || (5'd28/*MS*/==-11'd539+xpc10nz) || (5'd28/*MS*/==
              -11'd537+xpc10nz) || (5'd28/*MS*/==-11'd534+xpc10nz) || (5'd28/*MS*/==-11'd532+xpc10nz) || (5'd28/*MS*/==-11'd528+xpc10nz
              ) || (5'd28/*MS*/==-10'd503+xpc10nz) || (5'd28/*MS*/==-10'd502+xpc10nz) || (5'd28/*MS*/==-10'd472+xpc10nz) || (5'd28/*MS*/==
              -10'd407+xpc10nz) || (5'd28/*MS*/==-10'd342+xpc10nz) || (5'd28/*MS*/==-10'd341+xpc10nz) || (5'd28/*MS*/==-10'd340+xpc10nz
              ) || (5'd28/*MS*/==-10'd338+xpc10nz) || (5'd28/*MS*/==-10'd335+xpc10nz) || (5'd28/*MS*/==-10'd334+xpc10nz) || (5'd28/*MS*/==
              -10'd330+xpc10nz) || (5'd28/*MS*/==-10'd329+xpc10nz) || (5'd28/*MS*/==-10'd327+xpc10nz) || (5'd28/*MS*/==-10'd324+xpc10nz
              ) || (5'd28/*MS*/==-10'd323+xpc10nz) || (5'd28/*MS*/==-10'd322+xpc10nz) || (5'd28/*MS*/==-10'd321+xpc10nz) || (5'd28/*MS*/==
              -10'd320+xpc10nz) || (5'd28/*MS*/==-10'd319+xpc10nz) || (5'd28/*MS*/==-10'd318+xpc10nz) || (5'd28/*MS*/==-10'd314+xpc10nz
              ) || (5'd28/*MS*/==-10'd289+xpc10nz) || (5'd28/*MS*/==-10'd287+xpc10nz) || (5'd28/*MS*/==-10'd285+xpc10nz) || (5'd28/*MS*/==
              -10'd284+xpc10nz) || (5'd28/*MS*/==-10'd259+xpc10nz) || (5'd28/*MS*/==-10'd258+xpc10nz) || (5'd28/*MS*/==-10'd257+xpc10nz
              ) || (5'd28/*MS*/==-9'd255+xpc10nz) || (5'd28/*MS*/==-9'd254+xpc10nz) || (5'd28/*MS*/==-9'd253+xpc10nz) || (5'd28/*MS*/==
              -9'd252+xpc10nz) || (5'd28/*MS*/==-9'd251+xpc10nz) || (5'd28/*MS*/==-9'd250+xpc10nz) || (5'd28/*MS*/==-9'd249+xpc10nz) || 
              (5'd28/*MS*/==-9'd248+xpc10nz) || (5'd28/*MS*/==-9'd247+xpc10nz) || (5'd28/*MS*/==-9'd246+xpc10nz) || (5'd28/*MS*/==-9'd245
              +xpc10nz) || (5'd28/*MS*/==-9'd244+xpc10nz) || (5'd28/*MS*/==-9'd242+xpc10nz) || (5'd28/*MS*/==-9'd241+xpc10nz) || (5'd28
              /*MS*/==-9'd239+xpc10nz) || (5'd28/*MS*/==-9'd238+xpc10nz) || (5'd28/*MS*/==-9'd236+xpc10nz) || (5'd28/*MS*/==-9'd171+xpc10nz
              ) || (5'd28/*MS*/==-8'd106+xpc10nz) || (5'd28/*MS*/==-8'd105+xpc10nz) || (5'd28/*MS*/==-8'd104+xpc10nz) || (5'd28/*MS*/==
              -8'd103+xpc10nz) || (5'd28/*MS*/==-8'd102+xpc10nz) || (5'd28/*MS*/==-8'd101+xpc10nz) || (5'd28/*MS*/==-8'd100+xpc10nz) || 
              (5'd28/*MS*/==-8'd99+xpc10nz) || (5'd28/*MS*/==-8'd98+xpc10nz) || (5'd28/*MS*/==-8'd97+xpc10nz) || (5'd28/*MS*/==-8'd96
              +xpc10nz) || (5'd28/*MS*/==-8'd95+xpc10nz) || (5'd28/*MS*/==-8'd94+xpc10nz) || (5'd28/*MS*/==-8'd93+xpc10nz) || (5'd28/*MS*/==
              -8'd92+xpc10nz) || (5'd28/*MS*/==-8'd91+xpc10nz) || (5'd28/*MS*/==-8'd90+xpc10nz) || (5'd28/*MS*/==-8'd89+xpc10nz) || (5'd28
              /*MS*/==-8'd88+xpc10nz) || (5'd28/*MS*/==-8'd87+xpc10nz) || (5'd28/*MS*/==-8'd86+xpc10nz) || (5'd28/*MS*/==-8'd85+xpc10nz
              ) || (5'd28/*MS*/==-8'd84+xpc10nz) || (5'd28/*MS*/==-8'd83+xpc10nz) || (5'd28/*MS*/==-8'd82+xpc10nz) || (5'd28/*MS*/==-8'd65
              +xpc10nz) || (5'd28/*MS*/==-8'd64+xpc10nz) || (5'd28/*MS*/==-7'd59+xpc10nz) || (5'd28/*MS*/==-7'd50+xpc10nz) || (5'd28/*MS*/==
              -7'd37+xpc10nz) || (5'd28/*MS*/==-6'd20+xpc10nz) || (5'd28/*MS*/==-6'd19+xpc10nz) || (5'd28/*MS*/==-6'd18+xpc10nz) || (5'd28
              /*MS*/==-6'd17+xpc10nz) || (5'd28/*MS*/==-6'd16+xpc10nz) || (5'd28/*MS*/==-5'd15+xpc10nz) || (5'd28/*MS*/==-5'd14+xpc10nz
              ) || (5'd28/*MS*/==-5'd13+xpc10nz) || (5'd28/*MS*/==-5'd12+xpc10nz) || (5'd28/*MS*/==-5'd11+xpc10nz) || (5'd28/*MS*/==-5'd10
              +xpc10nz) || (5'd28/*MS*/==-5'd9+xpc10nz) || (5'd28/*MS*/==-5'd8+xpc10nz) || (5'd28/*MS*/==-4'd7+xpc10nz) || (5'd28/*MS*/==
              -4'd6+xpc10nz) || (5'd28/*MS*/==-4'd5+xpc10nz) || (5'd28/*MS*/==-4'd4+xpc10nz) || (5'd28/*MS*/==-3'd3+xpc10nz) || (5'd28
              /*MS*/==-3'd2+xpc10nz) || (5'd28/*MS*/==-2'd1+xpc10nz) || (xpc10nz==5'd28/*US*/)) && !xpc10_clear && !xpc10_stall;

               xpc10_trk27 <= ((5'd27/*MS*/==-11'd609+xpc10nz) || (5'd27/*MS*/==-11'd599+xpc10nz) || (5'd27/*MS*/==-11'd588+xpc10nz) || 
              (5'd27/*MS*/==-11'd576+xpc10nz) || (5'd27/*MS*/==-11'd571+xpc10nz) || (5'd27/*MS*/==-11'd565+xpc10nz) || (5'd27/*MS*/==
              -11'd558+xpc10nz) || (5'd27/*MS*/==-11'd550+xpc10nz) || (5'd27/*MS*/==-11'd549+xpc10nz) || (5'd27/*MS*/==-11'd547+xpc10nz
              ) || (5'd27/*MS*/==-11'd544+xpc10nz) || (5'd27/*MS*/==-11'd540+xpc10nz) || (5'd27/*MS*/==-11'd539+xpc10nz) || (5'd27/*MS*/==
              -11'd537+xpc10nz) || (5'd27/*MS*/==-11'd534+xpc10nz) || (5'd27/*MS*/==-11'd532+xpc10nz) || (5'd27/*MS*/==-11'd528+xpc10nz
              ) || (5'd27/*MS*/==-10'd503+xpc10nz) || (5'd27/*MS*/==-10'd502+xpc10nz) || (5'd27/*MS*/==-10'd472+xpc10nz) || (5'd27/*MS*/==
              -10'd407+xpc10nz) || (5'd27/*MS*/==-10'd342+xpc10nz) || (5'd27/*MS*/==-10'd341+xpc10nz) || (5'd27/*MS*/==-10'd340+xpc10nz
              ) || (5'd27/*MS*/==-10'd338+xpc10nz) || (5'd27/*MS*/==-10'd335+xpc10nz) || (5'd27/*MS*/==-10'd334+xpc10nz) || (5'd27/*MS*/==
              -10'd330+xpc10nz) || (5'd27/*MS*/==-10'd329+xpc10nz) || (5'd27/*MS*/==-10'd327+xpc10nz) || (5'd27/*MS*/==-10'd324+xpc10nz
              ) || (5'd27/*MS*/==-10'd323+xpc10nz) || (5'd27/*MS*/==-10'd322+xpc10nz) || (5'd27/*MS*/==-10'd321+xpc10nz) || (5'd27/*MS*/==
              -10'd320+xpc10nz) || (5'd27/*MS*/==-10'd319+xpc10nz) || (5'd27/*MS*/==-10'd318+xpc10nz) || (5'd27/*MS*/==-10'd314+xpc10nz
              ) || (5'd27/*MS*/==-10'd289+xpc10nz) || (5'd27/*MS*/==-10'd287+xpc10nz) || (5'd27/*MS*/==-10'd285+xpc10nz) || (5'd27/*MS*/==
              -10'd284+xpc10nz) || (5'd27/*MS*/==-10'd259+xpc10nz) || (5'd27/*MS*/==-10'd258+xpc10nz) || (5'd27/*MS*/==-10'd257+xpc10nz
              ) || (5'd27/*MS*/==-9'd255+xpc10nz) || (5'd27/*MS*/==-9'd254+xpc10nz) || (5'd27/*MS*/==-9'd253+xpc10nz) || (5'd27/*MS*/==
              -9'd252+xpc10nz) || (5'd27/*MS*/==-9'd251+xpc10nz) || (5'd27/*MS*/==-9'd250+xpc10nz) || (5'd27/*MS*/==-9'd249+xpc10nz) || 
              (5'd27/*MS*/==-9'd248+xpc10nz) || (5'd27/*MS*/==-9'd247+xpc10nz) || (5'd27/*MS*/==-9'd246+xpc10nz) || (5'd27/*MS*/==-9'd245
              +xpc10nz) || (5'd27/*MS*/==-9'd244+xpc10nz) || (5'd27/*MS*/==-9'd242+xpc10nz) || (5'd27/*MS*/==-9'd241+xpc10nz) || (5'd27
              /*MS*/==-9'd239+xpc10nz) || (5'd27/*MS*/==-9'd238+xpc10nz) || (5'd27/*MS*/==-9'd236+xpc10nz) || (5'd27/*MS*/==-9'd171+xpc10nz
              ) || (5'd27/*MS*/==-8'd106+xpc10nz) || (5'd27/*MS*/==-8'd105+xpc10nz) || (5'd27/*MS*/==-8'd104+xpc10nz) || (5'd27/*MS*/==
              -8'd103+xpc10nz) || (5'd27/*MS*/==-8'd102+xpc10nz) || (5'd27/*MS*/==-8'd101+xpc10nz) || (5'd27/*MS*/==-8'd100+xpc10nz) || 
              (5'd27/*MS*/==-8'd99+xpc10nz) || (5'd27/*MS*/==-8'd98+xpc10nz) || (5'd27/*MS*/==-8'd97+xpc10nz) || (5'd27/*MS*/==-8'd96
              +xpc10nz) || (5'd27/*MS*/==-8'd95+xpc10nz) || (5'd27/*MS*/==-8'd94+xpc10nz) || (5'd27/*MS*/==-8'd93+xpc10nz) || (5'd27/*MS*/==
              -8'd92+xpc10nz) || (5'd27/*MS*/==-8'd91+xpc10nz) || (5'd27/*MS*/==-8'd90+xpc10nz) || (5'd27/*MS*/==-8'd89+xpc10nz) || (5'd27
              /*MS*/==-8'd88+xpc10nz) || (5'd27/*MS*/==-8'd87+xpc10nz) || (5'd27/*MS*/==-8'd86+xpc10nz) || (5'd27/*MS*/==-8'd85+xpc10nz
              ) || (5'd27/*MS*/==-8'd84+xpc10nz) || (5'd27/*MS*/==-8'd83+xpc10nz) || (5'd27/*MS*/==-8'd82+xpc10nz) || (5'd27/*MS*/==-8'd65
              +xpc10nz) || (5'd27/*MS*/==-8'd64+xpc10nz) || (5'd27/*MS*/==-7'd59+xpc10nz) || (5'd27/*MS*/==-7'd50+xpc10nz) || (5'd27/*MS*/==
              -7'd37+xpc10nz) || (5'd27/*MS*/==-6'd20+xpc10nz) || (5'd27/*MS*/==-6'd19+xpc10nz) || (5'd27/*MS*/==-6'd18+xpc10nz) || (5'd27
              /*MS*/==-6'd17+xpc10nz) || (5'd27/*MS*/==-6'd16+xpc10nz) || (5'd27/*MS*/==-5'd15+xpc10nz) || (5'd27/*MS*/==-5'd14+xpc10nz
              ) || (5'd27/*MS*/==-5'd13+xpc10nz) || (5'd27/*MS*/==-5'd12+xpc10nz) || (5'd27/*MS*/==-5'd11+xpc10nz) || (5'd27/*MS*/==-5'd10
              +xpc10nz) || (5'd27/*MS*/==-5'd9+xpc10nz) || (5'd27/*MS*/==-5'd8+xpc10nz) || (5'd27/*MS*/==-4'd7+xpc10nz) || (5'd27/*MS*/==
              -4'd6+xpc10nz) || (5'd27/*MS*/==-4'd5+xpc10nz) || (5'd27/*MS*/==-4'd4+xpc10nz) || (5'd27/*MS*/==-3'd3+xpc10nz) || (5'd27
              /*MS*/==-3'd2+xpc10nz) || (5'd27/*MS*/==-2'd1+xpc10nz) || (xpc10nz==5'd27/*US*/)) && !xpc10_clear && !xpc10_stall;

               xpc10_trk26 <= ((5'd26/*MS*/==-11'd609+xpc10nz) || (5'd26/*MS*/==-11'd599+xpc10nz) || (5'd26/*MS*/==-11'd588+xpc10nz) || 
              (5'd26/*MS*/==-11'd576+xpc10nz) || (5'd26/*MS*/==-11'd571+xpc10nz) || (5'd26/*MS*/==-11'd565+xpc10nz) || (5'd26/*MS*/==
              -11'd558+xpc10nz) || (5'd26/*MS*/==-11'd550+xpc10nz) || (5'd26/*MS*/==-11'd549+xpc10nz) || (5'd26/*MS*/==-11'd547+xpc10nz
              ) || (5'd26/*MS*/==-11'd544+xpc10nz) || (5'd26/*MS*/==-11'd540+xpc10nz) || (5'd26/*MS*/==-11'd539+xpc10nz) || (5'd26/*MS*/==
              -11'd537+xpc10nz) || (5'd26/*MS*/==-11'd534+xpc10nz) || (5'd26/*MS*/==-11'd532+xpc10nz) || (5'd26/*MS*/==-11'd528+xpc10nz
              ) || (5'd26/*MS*/==-10'd503+xpc10nz) || (5'd26/*MS*/==-10'd502+xpc10nz) || (5'd26/*MS*/==-10'd472+xpc10nz) || (5'd26/*MS*/==
              -10'd407+xpc10nz) || (5'd26/*MS*/==-10'd342+xpc10nz) || (5'd26/*MS*/==-10'd341+xpc10nz) || (5'd26/*MS*/==-10'd340+xpc10nz
              ) || (5'd26/*MS*/==-10'd338+xpc10nz) || (5'd26/*MS*/==-10'd335+xpc10nz) || (5'd26/*MS*/==-10'd334+xpc10nz) || (5'd26/*MS*/==
              -10'd330+xpc10nz) || (5'd26/*MS*/==-10'd329+xpc10nz) || (5'd26/*MS*/==-10'd327+xpc10nz) || (5'd26/*MS*/==-10'd324+xpc10nz
              ) || (5'd26/*MS*/==-10'd323+xpc10nz) || (5'd26/*MS*/==-10'd322+xpc10nz) || (5'd26/*MS*/==-10'd321+xpc10nz) || (5'd26/*MS*/==
              -10'd320+xpc10nz) || (5'd26/*MS*/==-10'd319+xpc10nz) || (5'd26/*MS*/==-10'd318+xpc10nz) || (5'd26/*MS*/==-10'd314+xpc10nz
              ) || (5'd26/*MS*/==-10'd289+xpc10nz) || (5'd26/*MS*/==-10'd287+xpc10nz) || (5'd26/*MS*/==-10'd285+xpc10nz) || (5'd26/*MS*/==
              -10'd284+xpc10nz) || (5'd26/*MS*/==-10'd259+xpc10nz) || (5'd26/*MS*/==-10'd258+xpc10nz) || (5'd26/*MS*/==-10'd257+xpc10nz
              ) || (5'd26/*MS*/==-9'd255+xpc10nz) || (5'd26/*MS*/==-9'd254+xpc10nz) || (5'd26/*MS*/==-9'd253+xpc10nz) || (5'd26/*MS*/==
              -9'd252+xpc10nz) || (5'd26/*MS*/==-9'd251+xpc10nz) || (5'd26/*MS*/==-9'd250+xpc10nz) || (5'd26/*MS*/==-9'd249+xpc10nz) || 
              (5'd26/*MS*/==-9'd248+xpc10nz) || (5'd26/*MS*/==-9'd247+xpc10nz) || (5'd26/*MS*/==-9'd246+xpc10nz) || (5'd26/*MS*/==-9'd245
              +xpc10nz) || (5'd26/*MS*/==-9'd244+xpc10nz) || (5'd26/*MS*/==-9'd242+xpc10nz) || (5'd26/*MS*/==-9'd241+xpc10nz) || (5'd26
              /*MS*/==-9'd239+xpc10nz) || (5'd26/*MS*/==-9'd238+xpc10nz) || (5'd26/*MS*/==-9'd236+xpc10nz) || (5'd26/*MS*/==-9'd171+xpc10nz
              ) || (5'd26/*MS*/==-8'd106+xpc10nz) || (5'd26/*MS*/==-8'd105+xpc10nz) || (5'd26/*MS*/==-8'd104+xpc10nz) || (5'd26/*MS*/==
              -8'd103+xpc10nz) || (5'd26/*MS*/==-8'd102+xpc10nz) || (5'd26/*MS*/==-8'd101+xpc10nz) || (5'd26/*MS*/==-8'd100+xpc10nz) || 
              (5'd26/*MS*/==-8'd99+xpc10nz) || (5'd26/*MS*/==-8'd98+xpc10nz) || (5'd26/*MS*/==-8'd97+xpc10nz) || (5'd26/*MS*/==-8'd96
              +xpc10nz) || (5'd26/*MS*/==-8'd95+xpc10nz) || (5'd26/*MS*/==-8'd94+xpc10nz) || (5'd26/*MS*/==-8'd93+xpc10nz) || (5'd26/*MS*/==
              -8'd92+xpc10nz) || (5'd26/*MS*/==-8'd91+xpc10nz) || (5'd26/*MS*/==-8'd90+xpc10nz) || (5'd26/*MS*/==-8'd89+xpc10nz) || (5'd26
              /*MS*/==-8'd88+xpc10nz) || (5'd26/*MS*/==-8'd87+xpc10nz) || (5'd26/*MS*/==-8'd86+xpc10nz) || (5'd26/*MS*/==-8'd85+xpc10nz
              ) || (5'd26/*MS*/==-8'd84+xpc10nz) || (5'd26/*MS*/==-8'd83+xpc10nz) || (5'd26/*MS*/==-8'd82+xpc10nz) || (5'd26/*MS*/==-8'd65
              +xpc10nz) || (5'd26/*MS*/==-8'd64+xpc10nz) || (5'd26/*MS*/==-7'd59+xpc10nz) || (5'd26/*MS*/==-7'd50+xpc10nz) || (5'd26/*MS*/==
              -7'd37+xpc10nz) || (5'd26/*MS*/==-6'd20+xpc10nz) || (5'd26/*MS*/==-6'd19+xpc10nz) || (5'd26/*MS*/==-6'd18+xpc10nz) || (5'd26
              /*MS*/==-6'd17+xpc10nz) || (5'd26/*MS*/==-6'd16+xpc10nz) || (5'd26/*MS*/==-5'd15+xpc10nz) || (5'd26/*MS*/==-5'd14+xpc10nz
              ) || (5'd26/*MS*/==-5'd13+xpc10nz) || (5'd26/*MS*/==-5'd12+xpc10nz) || (5'd26/*MS*/==-5'd11+xpc10nz) || (5'd26/*MS*/==-5'd10
              +xpc10nz) || (5'd26/*MS*/==-5'd9+xpc10nz) || (5'd26/*MS*/==-5'd8+xpc10nz) || (5'd26/*MS*/==-4'd7+xpc10nz) || (5'd26/*MS*/==
              -4'd6+xpc10nz) || (5'd26/*MS*/==-4'd5+xpc10nz) || (5'd26/*MS*/==-4'd4+xpc10nz) || (5'd26/*MS*/==-3'd3+xpc10nz) || (5'd26
              /*MS*/==-3'd2+xpc10nz) || (5'd26/*MS*/==-2'd1+xpc10nz) || (xpc10nz==5'd26/*US*/)) && !xpc10_clear && !xpc10_stall;

               xpc10_trk25 <= ((5'd25/*MS*/==-11'd609+xpc10nz) || (5'd25/*MS*/==-11'd599+xpc10nz) || (5'd25/*MS*/==-11'd588+xpc10nz) || 
              (5'd25/*MS*/==-11'd576+xpc10nz) || (5'd25/*MS*/==-11'd571+xpc10nz) || (5'd25/*MS*/==-11'd565+xpc10nz) || (5'd25/*MS*/==
              -11'd558+xpc10nz) || (5'd25/*MS*/==-11'd550+xpc10nz) || (5'd25/*MS*/==-11'd549+xpc10nz) || (5'd25/*MS*/==-11'd547+xpc10nz
              ) || (5'd25/*MS*/==-11'd544+xpc10nz) || (5'd25/*MS*/==-11'd540+xpc10nz) || (5'd25/*MS*/==-11'd539+xpc10nz) || (5'd25/*MS*/==
              -11'd537+xpc10nz) || (5'd25/*MS*/==-11'd534+xpc10nz) || (5'd25/*MS*/==-11'd532+xpc10nz) || (5'd25/*MS*/==-11'd528+xpc10nz
              ) || (5'd25/*MS*/==-10'd503+xpc10nz) || (5'd25/*MS*/==-10'd502+xpc10nz) || (5'd25/*MS*/==-10'd472+xpc10nz) || (5'd25/*MS*/==
              -10'd407+xpc10nz) || (5'd25/*MS*/==-10'd342+xpc10nz) || (5'd25/*MS*/==-10'd341+xpc10nz) || (5'd25/*MS*/==-10'd340+xpc10nz
              ) || (5'd25/*MS*/==-10'd338+xpc10nz) || (5'd25/*MS*/==-10'd335+xpc10nz) || (5'd25/*MS*/==-10'd334+xpc10nz) || (5'd25/*MS*/==
              -10'd330+xpc10nz) || (5'd25/*MS*/==-10'd329+xpc10nz) || (5'd25/*MS*/==-10'd327+xpc10nz) || (5'd25/*MS*/==-10'd324+xpc10nz
              ) || (5'd25/*MS*/==-10'd323+xpc10nz) || (5'd25/*MS*/==-10'd322+xpc10nz) || (5'd25/*MS*/==-10'd321+xpc10nz) || (5'd25/*MS*/==
              -10'd320+xpc10nz) || (5'd25/*MS*/==-10'd319+xpc10nz) || (5'd25/*MS*/==-10'd318+xpc10nz) || (5'd25/*MS*/==-10'd314+xpc10nz
              ) || (5'd25/*MS*/==-10'd289+xpc10nz) || (5'd25/*MS*/==-10'd287+xpc10nz) || (5'd25/*MS*/==-10'd285+xpc10nz) || (5'd25/*MS*/==
              -10'd284+xpc10nz) || (5'd25/*MS*/==-10'd259+xpc10nz) || (5'd25/*MS*/==-10'd258+xpc10nz) || (5'd25/*MS*/==-10'd257+xpc10nz
              ) || (5'd25/*MS*/==-9'd255+xpc10nz) || (5'd25/*MS*/==-9'd254+xpc10nz) || (5'd25/*MS*/==-9'd253+xpc10nz) || (5'd25/*MS*/==
              -9'd252+xpc10nz) || (5'd25/*MS*/==-9'd251+xpc10nz) || (5'd25/*MS*/==-9'd250+xpc10nz) || (5'd25/*MS*/==-9'd249+xpc10nz) || 
              (5'd25/*MS*/==-9'd248+xpc10nz) || (5'd25/*MS*/==-9'd247+xpc10nz) || (5'd25/*MS*/==-9'd246+xpc10nz) || (5'd25/*MS*/==-9'd245
              +xpc10nz) || (5'd25/*MS*/==-9'd244+xpc10nz) || (5'd25/*MS*/==-9'd242+xpc10nz) || (5'd25/*MS*/==-9'd241+xpc10nz) || (5'd25
              /*MS*/==-9'd239+xpc10nz) || (5'd25/*MS*/==-9'd238+xpc10nz) || (5'd25/*MS*/==-9'd236+xpc10nz) || (5'd25/*MS*/==-9'd171+xpc10nz
              ) || (5'd25/*MS*/==-8'd106+xpc10nz) || (5'd25/*MS*/==-8'd105+xpc10nz) || (5'd25/*MS*/==-8'd104+xpc10nz) || (5'd25/*MS*/==
              -8'd103+xpc10nz) || (5'd25/*MS*/==-8'd102+xpc10nz) || (5'd25/*MS*/==-8'd101+xpc10nz) || (5'd25/*MS*/==-8'd100+xpc10nz) || 
              (5'd25/*MS*/==-8'd99+xpc10nz) || (5'd25/*MS*/==-8'd98+xpc10nz) || (5'd25/*MS*/==-8'd97+xpc10nz) || (5'd25/*MS*/==-8'd96
              +xpc10nz) || (5'd25/*MS*/==-8'd95+xpc10nz) || (5'd25/*MS*/==-8'd94+xpc10nz) || (5'd25/*MS*/==-8'd93+xpc10nz) || (5'd25/*MS*/==
              -8'd92+xpc10nz) || (5'd25/*MS*/==-8'd91+xpc10nz) || (5'd25/*MS*/==-8'd90+xpc10nz) || (5'd25/*MS*/==-8'd89+xpc10nz) || (5'd25
              /*MS*/==-8'd88+xpc10nz) || (5'd25/*MS*/==-8'd87+xpc10nz) || (5'd25/*MS*/==-8'd86+xpc10nz) || (5'd25/*MS*/==-8'd85+xpc10nz
              ) || (5'd25/*MS*/==-8'd84+xpc10nz) || (5'd25/*MS*/==-8'd83+xpc10nz) || (5'd25/*MS*/==-8'd82+xpc10nz) || (5'd25/*MS*/==-8'd65
              +xpc10nz) || (5'd25/*MS*/==-8'd64+xpc10nz) || (5'd25/*MS*/==-7'd59+xpc10nz) || (5'd25/*MS*/==-7'd50+xpc10nz) || (5'd25/*MS*/==
              -7'd37+xpc10nz) || (5'd25/*MS*/==-6'd20+xpc10nz) || (5'd25/*MS*/==-6'd19+xpc10nz) || (5'd25/*MS*/==-6'd18+xpc10nz) || (5'd25
              /*MS*/==-6'd17+xpc10nz) || (5'd25/*MS*/==-6'd16+xpc10nz) || (5'd25/*MS*/==-5'd15+xpc10nz) || (5'd25/*MS*/==-5'd14+xpc10nz
              ) || (5'd25/*MS*/==-5'd13+xpc10nz) || (5'd25/*MS*/==-5'd12+xpc10nz) || (5'd25/*MS*/==-5'd11+xpc10nz) || (5'd25/*MS*/==-5'd10
              +xpc10nz) || (5'd25/*MS*/==-5'd9+xpc10nz) || (5'd25/*MS*/==-5'd8+xpc10nz) || (5'd25/*MS*/==-4'd7+xpc10nz) || (5'd25/*MS*/==
              -4'd6+xpc10nz) || (5'd25/*MS*/==-4'd5+xpc10nz) || (5'd25/*MS*/==-4'd4+xpc10nz) || (5'd25/*MS*/==-3'd3+xpc10nz) || (5'd25
              /*MS*/==-3'd2+xpc10nz) || (5'd25/*MS*/==-2'd1+xpc10nz) || (xpc10nz==5'd25/*US*/)) && !xpc10_clear && !xpc10_stall;

               xpc10_trk24 <= ((5'd24/*MS*/==-11'd609+xpc10nz) || (5'd24/*MS*/==-11'd599+xpc10nz) || (5'd24/*MS*/==-11'd588+xpc10nz) || 
              (5'd24/*MS*/==-11'd576+xpc10nz) || (5'd24/*MS*/==-11'd571+xpc10nz) || (5'd24/*MS*/==-11'd565+xpc10nz) || (5'd24/*MS*/==
              -11'd558+xpc10nz) || (5'd24/*MS*/==-11'd550+xpc10nz) || (5'd24/*MS*/==-11'd549+xpc10nz) || (5'd24/*MS*/==-11'd547+xpc10nz
              ) || (5'd24/*MS*/==-11'd544+xpc10nz) || (5'd24/*MS*/==-11'd540+xpc10nz) || (5'd24/*MS*/==-11'd539+xpc10nz) || (5'd24/*MS*/==
              -11'd537+xpc10nz) || (5'd24/*MS*/==-11'd534+xpc10nz) || (5'd24/*MS*/==-11'd532+xpc10nz) || (5'd24/*MS*/==-11'd528+xpc10nz
              ) || (5'd24/*MS*/==-10'd503+xpc10nz) || (5'd24/*MS*/==-10'd502+xpc10nz) || (5'd24/*MS*/==-10'd472+xpc10nz) || (5'd24/*MS*/==
              -10'd407+xpc10nz) || (5'd24/*MS*/==-10'd342+xpc10nz) || (5'd24/*MS*/==-10'd341+xpc10nz) || (5'd24/*MS*/==-10'd340+xpc10nz
              ) || (5'd24/*MS*/==-10'd338+xpc10nz) || (5'd24/*MS*/==-10'd335+xpc10nz) || (5'd24/*MS*/==-10'd334+xpc10nz) || (5'd24/*MS*/==
              -10'd330+xpc10nz) || (5'd24/*MS*/==-10'd329+xpc10nz) || (5'd24/*MS*/==-10'd327+xpc10nz) || (5'd24/*MS*/==-10'd324+xpc10nz
              ) || (5'd24/*MS*/==-10'd323+xpc10nz) || (5'd24/*MS*/==-10'd322+xpc10nz) || (5'd24/*MS*/==-10'd321+xpc10nz) || (5'd24/*MS*/==
              -10'd320+xpc10nz) || (5'd24/*MS*/==-10'd319+xpc10nz) || (5'd24/*MS*/==-10'd318+xpc10nz) || (5'd24/*MS*/==-10'd314+xpc10nz
              ) || (5'd24/*MS*/==-10'd289+xpc10nz) || (5'd24/*MS*/==-10'd287+xpc10nz) || (5'd24/*MS*/==-10'd285+xpc10nz) || (5'd24/*MS*/==
              -10'd284+xpc10nz) || (5'd24/*MS*/==-10'd259+xpc10nz) || (5'd24/*MS*/==-10'd258+xpc10nz) || (5'd24/*MS*/==-10'd257+xpc10nz
              ) || (5'd24/*MS*/==-9'd255+xpc10nz) || (5'd24/*MS*/==-9'd254+xpc10nz) || (5'd24/*MS*/==-9'd253+xpc10nz) || (5'd24/*MS*/==
              -9'd252+xpc10nz) || (5'd24/*MS*/==-9'd251+xpc10nz) || (5'd24/*MS*/==-9'd250+xpc10nz) || (5'd24/*MS*/==-9'd249+xpc10nz) || 
              (5'd24/*MS*/==-9'd248+xpc10nz) || (5'd24/*MS*/==-9'd247+xpc10nz) || (5'd24/*MS*/==-9'd246+xpc10nz) || (5'd24/*MS*/==-9'd245
              +xpc10nz) || (5'd24/*MS*/==-9'd244+xpc10nz) || (5'd24/*MS*/==-9'd242+xpc10nz) || (5'd24/*MS*/==-9'd241+xpc10nz) || (5'd24
              /*MS*/==-9'd239+xpc10nz) || (5'd24/*MS*/==-9'd238+xpc10nz) || (5'd24/*MS*/==-9'd236+xpc10nz) || (5'd24/*MS*/==-9'd171+xpc10nz
              ) || (5'd24/*MS*/==-8'd106+xpc10nz) || (5'd24/*MS*/==-8'd105+xpc10nz) || (5'd24/*MS*/==-8'd104+xpc10nz) || (5'd24/*MS*/==
              -8'd103+xpc10nz) || (5'd24/*MS*/==-8'd102+xpc10nz) || (5'd24/*MS*/==-8'd101+xpc10nz) || (5'd24/*MS*/==-8'd100+xpc10nz) || 
              (5'd24/*MS*/==-8'd99+xpc10nz) || (5'd24/*MS*/==-8'd98+xpc10nz) || (5'd24/*MS*/==-8'd97+xpc10nz) || (5'd24/*MS*/==-8'd96
              +xpc10nz) || (5'd24/*MS*/==-8'd95+xpc10nz) || (5'd24/*MS*/==-8'd94+xpc10nz) || (5'd24/*MS*/==-8'd93+xpc10nz) || (5'd24/*MS*/==
              -8'd92+xpc10nz) || (5'd24/*MS*/==-8'd91+xpc10nz) || (5'd24/*MS*/==-8'd90+xpc10nz) || (5'd24/*MS*/==-8'd89+xpc10nz) || (5'd24
              /*MS*/==-8'd88+xpc10nz) || (5'd24/*MS*/==-8'd87+xpc10nz) || (5'd24/*MS*/==-8'd86+xpc10nz) || (5'd24/*MS*/==-8'd85+xpc10nz
              ) || (5'd24/*MS*/==-8'd84+xpc10nz) || (5'd24/*MS*/==-8'd83+xpc10nz) || (5'd24/*MS*/==-8'd82+xpc10nz) || (5'd24/*MS*/==-8'd65
              +xpc10nz) || (5'd24/*MS*/==-8'd64+xpc10nz) || (5'd24/*MS*/==-7'd59+xpc10nz) || (5'd24/*MS*/==-7'd50+xpc10nz) || (5'd24/*MS*/==
              -7'd37+xpc10nz) || (5'd24/*MS*/==-6'd20+xpc10nz) || (5'd24/*MS*/==-6'd19+xpc10nz) || (5'd24/*MS*/==-6'd18+xpc10nz) || (5'd24
              /*MS*/==-6'd17+xpc10nz) || (5'd24/*MS*/==-6'd16+xpc10nz) || (5'd24/*MS*/==-5'd15+xpc10nz) || (5'd24/*MS*/==-5'd14+xpc10nz
              ) || (5'd24/*MS*/==-5'd13+xpc10nz) || (5'd24/*MS*/==-5'd12+xpc10nz) || (5'd24/*MS*/==-5'd11+xpc10nz) || (5'd24/*MS*/==-5'd10
              +xpc10nz) || (5'd24/*MS*/==-5'd9+xpc10nz) || (5'd24/*MS*/==-5'd8+xpc10nz) || (5'd24/*MS*/==-4'd7+xpc10nz) || (5'd24/*MS*/==
              -4'd6+xpc10nz) || (5'd24/*MS*/==-4'd5+xpc10nz) || (5'd24/*MS*/==-4'd4+xpc10nz) || (5'd24/*MS*/==-3'd3+xpc10nz) || (5'd24
              /*MS*/==-3'd2+xpc10nz) || (5'd24/*MS*/==-2'd1+xpc10nz) || (xpc10nz==5'd24/*US*/)) && !xpc10_clear && !xpc10_stall;

               xpc10_trk23 <= ((5'd23/*MS*/==-11'd609+xpc10nz) || (5'd23/*MS*/==-11'd599+xpc10nz) || (5'd23/*MS*/==-11'd588+xpc10nz) || 
              (5'd23/*MS*/==-11'd576+xpc10nz) || (5'd23/*MS*/==-11'd571+xpc10nz) || (5'd23/*MS*/==-11'd565+xpc10nz) || (5'd23/*MS*/==
              -11'd558+xpc10nz) || (5'd23/*MS*/==-11'd550+xpc10nz) || (5'd23/*MS*/==-11'd549+xpc10nz) || (5'd23/*MS*/==-11'd547+xpc10nz
              ) || (5'd23/*MS*/==-11'd544+xpc10nz) || (5'd23/*MS*/==-11'd540+xpc10nz) || (5'd23/*MS*/==-11'd539+xpc10nz) || (5'd23/*MS*/==
              -11'd537+xpc10nz) || (5'd23/*MS*/==-11'd534+xpc10nz) || (5'd23/*MS*/==-11'd532+xpc10nz) || (5'd23/*MS*/==-11'd528+xpc10nz
              ) || (5'd23/*MS*/==-10'd503+xpc10nz) || (5'd23/*MS*/==-10'd502+xpc10nz) || (5'd23/*MS*/==-10'd472+xpc10nz) || (5'd23/*MS*/==
              -10'd407+xpc10nz) || (5'd23/*MS*/==-10'd342+xpc10nz) || (5'd23/*MS*/==-10'd341+xpc10nz) || (5'd23/*MS*/==-10'd340+xpc10nz
              ) || (5'd23/*MS*/==-10'd338+xpc10nz) || (5'd23/*MS*/==-10'd335+xpc10nz) || (5'd23/*MS*/==-10'd334+xpc10nz) || (5'd23/*MS*/==
              -10'd330+xpc10nz) || (5'd23/*MS*/==-10'd329+xpc10nz) || (5'd23/*MS*/==-10'd327+xpc10nz) || (5'd23/*MS*/==-10'd324+xpc10nz
              ) || (5'd23/*MS*/==-10'd323+xpc10nz) || (5'd23/*MS*/==-10'd322+xpc10nz) || (5'd23/*MS*/==-10'd321+xpc10nz) || (5'd23/*MS*/==
              -10'd320+xpc10nz) || (5'd23/*MS*/==-10'd319+xpc10nz) || (5'd23/*MS*/==-10'd318+xpc10nz) || (5'd23/*MS*/==-10'd314+xpc10nz
              ) || (5'd23/*MS*/==-10'd289+xpc10nz) || (5'd23/*MS*/==-10'd287+xpc10nz) || (5'd23/*MS*/==-10'd285+xpc10nz) || (5'd23/*MS*/==
              -10'd284+xpc10nz) || (5'd23/*MS*/==-10'd259+xpc10nz) || (5'd23/*MS*/==-10'd258+xpc10nz) || (5'd23/*MS*/==-10'd257+xpc10nz
              ) || (5'd23/*MS*/==-9'd255+xpc10nz) || (5'd23/*MS*/==-9'd254+xpc10nz) || (5'd23/*MS*/==-9'd253+xpc10nz) || (5'd23/*MS*/==
              -9'd252+xpc10nz) || (5'd23/*MS*/==-9'd251+xpc10nz) || (5'd23/*MS*/==-9'd250+xpc10nz) || (5'd23/*MS*/==-9'd249+xpc10nz) || 
              (5'd23/*MS*/==-9'd248+xpc10nz) || (5'd23/*MS*/==-9'd247+xpc10nz) || (5'd23/*MS*/==-9'd246+xpc10nz) || (5'd23/*MS*/==-9'd245
              +xpc10nz) || (5'd23/*MS*/==-9'd244+xpc10nz) || (5'd23/*MS*/==-9'd242+xpc10nz) || (5'd23/*MS*/==-9'd241+xpc10nz) || (5'd23
              /*MS*/==-9'd239+xpc10nz) || (5'd23/*MS*/==-9'd238+xpc10nz) || (5'd23/*MS*/==-9'd236+xpc10nz) || (5'd23/*MS*/==-9'd171+xpc10nz
              ) || (5'd23/*MS*/==-8'd106+xpc10nz) || (5'd23/*MS*/==-8'd105+xpc10nz) || (5'd23/*MS*/==-8'd104+xpc10nz) || (5'd23/*MS*/==
              -8'd103+xpc10nz) || (5'd23/*MS*/==-8'd102+xpc10nz) || (5'd23/*MS*/==-8'd101+xpc10nz) || (5'd23/*MS*/==-8'd100+xpc10nz) || 
              (5'd23/*MS*/==-8'd99+xpc10nz) || (5'd23/*MS*/==-8'd98+xpc10nz) || (5'd23/*MS*/==-8'd97+xpc10nz) || (5'd23/*MS*/==-8'd96
              +xpc10nz) || (5'd23/*MS*/==-8'd95+xpc10nz) || (5'd23/*MS*/==-8'd94+xpc10nz) || (5'd23/*MS*/==-8'd93+xpc10nz) || (5'd23/*MS*/==
              -8'd92+xpc10nz) || (5'd23/*MS*/==-8'd91+xpc10nz) || (5'd23/*MS*/==-8'd90+xpc10nz) || (5'd23/*MS*/==-8'd89+xpc10nz) || (5'd23
              /*MS*/==-8'd88+xpc10nz) || (5'd23/*MS*/==-8'd87+xpc10nz) || (5'd23/*MS*/==-8'd86+xpc10nz) || (5'd23/*MS*/==-8'd85+xpc10nz
              ) || (5'd23/*MS*/==-8'd84+xpc10nz) || (5'd23/*MS*/==-8'd83+xpc10nz) || (5'd23/*MS*/==-8'd82+xpc10nz) || (5'd23/*MS*/==-8'd65
              +xpc10nz) || (5'd23/*MS*/==-8'd64+xpc10nz) || (5'd23/*MS*/==-7'd59+xpc10nz) || (5'd23/*MS*/==-7'd50+xpc10nz) || (5'd23/*MS*/==
              -7'd37+xpc10nz) || (5'd23/*MS*/==-6'd20+xpc10nz) || (5'd23/*MS*/==-6'd19+xpc10nz) || (5'd23/*MS*/==-6'd18+xpc10nz) || (5'd23
              /*MS*/==-6'd17+xpc10nz) || (5'd23/*MS*/==-6'd16+xpc10nz) || (5'd23/*MS*/==-5'd15+xpc10nz) || (5'd23/*MS*/==-5'd14+xpc10nz
              ) || (5'd23/*MS*/==-5'd13+xpc10nz) || (5'd23/*MS*/==-5'd12+xpc10nz) || (5'd23/*MS*/==-5'd11+xpc10nz) || (5'd23/*MS*/==-5'd10
              +xpc10nz) || (5'd23/*MS*/==-5'd9+xpc10nz) || (5'd23/*MS*/==-5'd8+xpc10nz) || (5'd23/*MS*/==-4'd7+xpc10nz) || (5'd23/*MS*/==
              -4'd6+xpc10nz) || (5'd23/*MS*/==-4'd5+xpc10nz) || (5'd23/*MS*/==-4'd4+xpc10nz) || (5'd23/*MS*/==-3'd3+xpc10nz) || (5'd23
              /*MS*/==-3'd2+xpc10nz) || (5'd23/*MS*/==-2'd1+xpc10nz) || (xpc10nz==5'd23/*US*/)) && !xpc10_clear && !xpc10_stall;

               xpc10_trk22 <= ((5'd22/*MS*/==-11'd609+xpc10nz) || (5'd22/*MS*/==-11'd599+xpc10nz) || (5'd22/*MS*/==-11'd588+xpc10nz) || 
              (5'd22/*MS*/==-11'd576+xpc10nz) || (5'd22/*MS*/==-11'd571+xpc10nz) || (5'd22/*MS*/==-11'd565+xpc10nz) || (5'd22/*MS*/==
              -11'd558+xpc10nz) || (5'd22/*MS*/==-11'd550+xpc10nz) || (5'd22/*MS*/==-11'd549+xpc10nz) || (5'd22/*MS*/==-11'd547+xpc10nz
              ) || (5'd22/*MS*/==-11'd544+xpc10nz) || (5'd22/*MS*/==-11'd540+xpc10nz) || (5'd22/*MS*/==-11'd539+xpc10nz) || (5'd22/*MS*/==
              -11'd537+xpc10nz) || (5'd22/*MS*/==-11'd534+xpc10nz) || (5'd22/*MS*/==-11'd532+xpc10nz) || (5'd22/*MS*/==-11'd528+xpc10nz
              ) || (5'd22/*MS*/==-10'd503+xpc10nz) || (5'd22/*MS*/==-10'd502+xpc10nz) || (5'd22/*MS*/==-10'd472+xpc10nz) || (5'd22/*MS*/==
              -10'd407+xpc10nz) || (5'd22/*MS*/==-10'd342+xpc10nz) || (5'd22/*MS*/==-10'd341+xpc10nz) || (5'd22/*MS*/==-10'd340+xpc10nz
              ) || (5'd22/*MS*/==-10'd338+xpc10nz) || (5'd22/*MS*/==-10'd335+xpc10nz) || (5'd22/*MS*/==-10'd334+xpc10nz) || (5'd22/*MS*/==
              -10'd330+xpc10nz) || (5'd22/*MS*/==-10'd329+xpc10nz) || (5'd22/*MS*/==-10'd327+xpc10nz) || (5'd22/*MS*/==-10'd324+xpc10nz
              ) || (5'd22/*MS*/==-10'd323+xpc10nz) || (5'd22/*MS*/==-10'd322+xpc10nz) || (5'd22/*MS*/==-10'd321+xpc10nz) || (5'd22/*MS*/==
              -10'd320+xpc10nz) || (5'd22/*MS*/==-10'd319+xpc10nz) || (5'd22/*MS*/==-10'd318+xpc10nz) || (5'd22/*MS*/==-10'd314+xpc10nz
              ) || (5'd22/*MS*/==-10'd289+xpc10nz) || (5'd22/*MS*/==-10'd287+xpc10nz) || (5'd22/*MS*/==-10'd285+xpc10nz) || (5'd22/*MS*/==
              -10'd284+xpc10nz) || (5'd22/*MS*/==-10'd259+xpc10nz) || (5'd22/*MS*/==-10'd258+xpc10nz) || (5'd22/*MS*/==-10'd257+xpc10nz
              ) || (5'd22/*MS*/==-9'd255+xpc10nz) || (5'd22/*MS*/==-9'd254+xpc10nz) || (5'd22/*MS*/==-9'd253+xpc10nz) || (5'd22/*MS*/==
              -9'd252+xpc10nz) || (5'd22/*MS*/==-9'd251+xpc10nz) || (5'd22/*MS*/==-9'd250+xpc10nz) || (5'd22/*MS*/==-9'd249+xpc10nz) || 
              (5'd22/*MS*/==-9'd248+xpc10nz) || (5'd22/*MS*/==-9'd247+xpc10nz) || (5'd22/*MS*/==-9'd246+xpc10nz) || (5'd22/*MS*/==-9'd245
              +xpc10nz) || (5'd22/*MS*/==-9'd244+xpc10nz) || (5'd22/*MS*/==-9'd242+xpc10nz) || (5'd22/*MS*/==-9'd241+xpc10nz) || (5'd22
              /*MS*/==-9'd239+xpc10nz) || (5'd22/*MS*/==-9'd238+xpc10nz) || (5'd22/*MS*/==-9'd236+xpc10nz) || (5'd22/*MS*/==-9'd171+xpc10nz
              ) || (5'd22/*MS*/==-8'd106+xpc10nz) || (5'd22/*MS*/==-8'd105+xpc10nz) || (5'd22/*MS*/==-8'd104+xpc10nz) || (5'd22/*MS*/==
              -8'd103+xpc10nz) || (5'd22/*MS*/==-8'd102+xpc10nz) || (5'd22/*MS*/==-8'd101+xpc10nz) || (5'd22/*MS*/==-8'd100+xpc10nz) || 
              (5'd22/*MS*/==-8'd99+xpc10nz) || (5'd22/*MS*/==-8'd98+xpc10nz) || (5'd22/*MS*/==-8'd97+xpc10nz) || (5'd22/*MS*/==-8'd96
              +xpc10nz) || (5'd22/*MS*/==-8'd95+xpc10nz) || (5'd22/*MS*/==-8'd94+xpc10nz) || (5'd22/*MS*/==-8'd93+xpc10nz) || (5'd22/*MS*/==
              -8'd92+xpc10nz) || (5'd22/*MS*/==-8'd91+xpc10nz) || (5'd22/*MS*/==-8'd90+xpc10nz) || (5'd22/*MS*/==-8'd89+xpc10nz) || (5'd22
              /*MS*/==-8'd88+xpc10nz) || (5'd22/*MS*/==-8'd87+xpc10nz) || (5'd22/*MS*/==-8'd86+xpc10nz) || (5'd22/*MS*/==-8'd85+xpc10nz
              ) || (5'd22/*MS*/==-8'd84+xpc10nz) || (5'd22/*MS*/==-8'd83+xpc10nz) || (5'd22/*MS*/==-8'd82+xpc10nz) || (5'd22/*MS*/==-8'd65
              +xpc10nz) || (5'd22/*MS*/==-8'd64+xpc10nz) || (5'd22/*MS*/==-7'd59+xpc10nz) || (5'd22/*MS*/==-7'd50+xpc10nz) || (5'd22/*MS*/==
              -7'd37+xpc10nz) || (5'd22/*MS*/==-6'd20+xpc10nz) || (5'd22/*MS*/==-6'd19+xpc10nz) || (5'd22/*MS*/==-6'd18+xpc10nz) || (5'd22
              /*MS*/==-6'd17+xpc10nz) || (5'd22/*MS*/==-6'd16+xpc10nz) || (5'd22/*MS*/==-5'd15+xpc10nz) || (5'd22/*MS*/==-5'd14+xpc10nz
              ) || (5'd22/*MS*/==-5'd13+xpc10nz) || (5'd22/*MS*/==-5'd12+xpc10nz) || (5'd22/*MS*/==-5'd11+xpc10nz) || (5'd22/*MS*/==-5'd10
              +xpc10nz) || (5'd22/*MS*/==-5'd9+xpc10nz) || (5'd22/*MS*/==-5'd8+xpc10nz) || (5'd22/*MS*/==-4'd7+xpc10nz) || (5'd22/*MS*/==
              -4'd6+xpc10nz) || (5'd22/*MS*/==-4'd5+xpc10nz) || (5'd22/*MS*/==-4'd4+xpc10nz) || (5'd22/*MS*/==-3'd3+xpc10nz) || (5'd22
              /*MS*/==-3'd2+xpc10nz) || (5'd22/*MS*/==-2'd1+xpc10nz) || (xpc10nz==5'd22/*US*/)) && !xpc10_clear && !xpc10_stall;

               xpc10_trk21 <= ((5'd21/*MS*/==-11'd609+xpc10nz) || (5'd21/*MS*/==-11'd599+xpc10nz) || (5'd21/*MS*/==-11'd588+xpc10nz) || 
              (5'd21/*MS*/==-11'd576+xpc10nz) || (5'd21/*MS*/==-11'd571+xpc10nz) || (5'd21/*MS*/==-11'd565+xpc10nz) || (5'd21/*MS*/==
              -11'd558+xpc10nz) || (5'd21/*MS*/==-11'd550+xpc10nz) || (5'd21/*MS*/==-11'd549+xpc10nz) || (5'd21/*MS*/==-11'd547+xpc10nz
              ) || (5'd21/*MS*/==-11'd544+xpc10nz) || (5'd21/*MS*/==-11'd540+xpc10nz) || (5'd21/*MS*/==-11'd539+xpc10nz) || (5'd21/*MS*/==
              -11'd537+xpc10nz) || (5'd21/*MS*/==-11'd534+xpc10nz) || (5'd21/*MS*/==-11'd532+xpc10nz) || (5'd21/*MS*/==-11'd528+xpc10nz
              ) || (5'd21/*MS*/==-10'd503+xpc10nz) || (5'd21/*MS*/==-10'd502+xpc10nz) || (5'd21/*MS*/==-10'd472+xpc10nz) || (5'd21/*MS*/==
              -10'd407+xpc10nz) || (5'd21/*MS*/==-10'd342+xpc10nz) || (5'd21/*MS*/==-10'd341+xpc10nz) || (5'd21/*MS*/==-10'd340+xpc10nz
              ) || (5'd21/*MS*/==-10'd338+xpc10nz) || (5'd21/*MS*/==-10'd335+xpc10nz) || (5'd21/*MS*/==-10'd334+xpc10nz) || (5'd21/*MS*/==
              -10'd330+xpc10nz) || (5'd21/*MS*/==-10'd329+xpc10nz) || (5'd21/*MS*/==-10'd327+xpc10nz) || (5'd21/*MS*/==-10'd324+xpc10nz
              ) || (5'd21/*MS*/==-10'd323+xpc10nz) || (5'd21/*MS*/==-10'd322+xpc10nz) || (5'd21/*MS*/==-10'd321+xpc10nz) || (5'd21/*MS*/==
              -10'd320+xpc10nz) || (5'd21/*MS*/==-10'd319+xpc10nz) || (5'd21/*MS*/==-10'd318+xpc10nz) || (5'd21/*MS*/==-10'd314+xpc10nz
              ) || (5'd21/*MS*/==-10'd289+xpc10nz) || (5'd21/*MS*/==-10'd287+xpc10nz) || (5'd21/*MS*/==-10'd285+xpc10nz) || (5'd21/*MS*/==
              -10'd284+xpc10nz) || (5'd21/*MS*/==-10'd259+xpc10nz) || (5'd21/*MS*/==-10'd258+xpc10nz) || (5'd21/*MS*/==-10'd257+xpc10nz
              ) || (5'd21/*MS*/==-9'd255+xpc10nz) || (5'd21/*MS*/==-9'd254+xpc10nz) || (5'd21/*MS*/==-9'd253+xpc10nz) || (5'd21/*MS*/==
              -9'd252+xpc10nz) || (5'd21/*MS*/==-9'd251+xpc10nz) || (5'd21/*MS*/==-9'd250+xpc10nz) || (5'd21/*MS*/==-9'd249+xpc10nz) || 
              (5'd21/*MS*/==-9'd248+xpc10nz) || (5'd21/*MS*/==-9'd247+xpc10nz) || (5'd21/*MS*/==-9'd246+xpc10nz) || (5'd21/*MS*/==-9'd245
              +xpc10nz) || (5'd21/*MS*/==-9'd244+xpc10nz) || (5'd21/*MS*/==-9'd242+xpc10nz) || (5'd21/*MS*/==-9'd241+xpc10nz) || (5'd21
              /*MS*/==-9'd239+xpc10nz) || (5'd21/*MS*/==-9'd238+xpc10nz) || (5'd21/*MS*/==-9'd236+xpc10nz) || (5'd21/*MS*/==-9'd171+xpc10nz
              ) || (5'd21/*MS*/==-8'd106+xpc10nz) || (5'd21/*MS*/==-8'd105+xpc10nz) || (5'd21/*MS*/==-8'd104+xpc10nz) || (5'd21/*MS*/==
              -8'd103+xpc10nz) || (5'd21/*MS*/==-8'd102+xpc10nz) || (5'd21/*MS*/==-8'd101+xpc10nz) || (5'd21/*MS*/==-8'd100+xpc10nz) || 
              (5'd21/*MS*/==-8'd99+xpc10nz) || (5'd21/*MS*/==-8'd98+xpc10nz) || (5'd21/*MS*/==-8'd97+xpc10nz) || (5'd21/*MS*/==-8'd96
              +xpc10nz) || (5'd21/*MS*/==-8'd95+xpc10nz) || (5'd21/*MS*/==-8'd94+xpc10nz) || (5'd21/*MS*/==-8'd93+xpc10nz) || (5'd21/*MS*/==
              -8'd92+xpc10nz) || (5'd21/*MS*/==-8'd91+xpc10nz) || (5'd21/*MS*/==-8'd90+xpc10nz) || (5'd21/*MS*/==-8'd89+xpc10nz) || (5'd21
              /*MS*/==-8'd88+xpc10nz) || (5'd21/*MS*/==-8'd87+xpc10nz) || (5'd21/*MS*/==-8'd86+xpc10nz) || (5'd21/*MS*/==-8'd85+xpc10nz
              ) || (5'd21/*MS*/==-8'd84+xpc10nz) || (5'd21/*MS*/==-8'd83+xpc10nz) || (5'd21/*MS*/==-8'd82+xpc10nz) || (5'd21/*MS*/==-8'd65
              +xpc10nz) || (5'd21/*MS*/==-8'd64+xpc10nz) || (5'd21/*MS*/==-7'd59+xpc10nz) || (5'd21/*MS*/==-7'd50+xpc10nz) || (5'd21/*MS*/==
              -7'd37+xpc10nz) || (5'd21/*MS*/==-6'd20+xpc10nz) || (5'd21/*MS*/==-6'd19+xpc10nz) || (5'd21/*MS*/==-6'd18+xpc10nz) || (5'd21
              /*MS*/==-6'd17+xpc10nz) || (5'd21/*MS*/==-6'd16+xpc10nz) || (5'd21/*MS*/==-5'd15+xpc10nz) || (5'd21/*MS*/==-5'd14+xpc10nz
              ) || (5'd21/*MS*/==-5'd13+xpc10nz) || (5'd21/*MS*/==-5'd12+xpc10nz) || (5'd21/*MS*/==-5'd11+xpc10nz) || (5'd21/*MS*/==-5'd10
              +xpc10nz) || (5'd21/*MS*/==-5'd9+xpc10nz) || (5'd21/*MS*/==-5'd8+xpc10nz) || (5'd21/*MS*/==-4'd7+xpc10nz) || (5'd21/*MS*/==
              -4'd6+xpc10nz) || (5'd21/*MS*/==-4'd5+xpc10nz) || (5'd21/*MS*/==-4'd4+xpc10nz) || (5'd21/*MS*/==-3'd3+xpc10nz) || (5'd21
              /*MS*/==-3'd2+xpc10nz) || (5'd21/*MS*/==-2'd1+xpc10nz) || (xpc10nz==5'd21/*US*/)) && !xpc10_clear && !xpc10_stall;

               xpc10_trk20 <= ((5'd20/*MS*/==-11'd609+xpc10nz) || (5'd20/*MS*/==-11'd599+xpc10nz) || (5'd20/*MS*/==-11'd588+xpc10nz) || 
              (5'd20/*MS*/==-11'd576+xpc10nz) || (5'd20/*MS*/==-11'd571+xpc10nz) || (5'd20/*MS*/==-11'd565+xpc10nz) || (5'd20/*MS*/==
              -11'd558+xpc10nz) || (5'd20/*MS*/==-11'd550+xpc10nz) || (5'd20/*MS*/==-11'd549+xpc10nz) || (5'd20/*MS*/==-11'd547+xpc10nz
              ) || (5'd20/*MS*/==-11'd544+xpc10nz) || (5'd20/*MS*/==-11'd540+xpc10nz) || (5'd20/*MS*/==-11'd539+xpc10nz) || (5'd20/*MS*/==
              -11'd537+xpc10nz) || (5'd20/*MS*/==-11'd534+xpc10nz) || (5'd20/*MS*/==-11'd532+xpc10nz) || (5'd20/*MS*/==-11'd528+xpc10nz
              ) || (5'd20/*MS*/==-10'd503+xpc10nz) || (5'd20/*MS*/==-10'd502+xpc10nz) || (5'd20/*MS*/==-10'd472+xpc10nz) || (5'd20/*MS*/==
              -10'd407+xpc10nz) || (5'd20/*MS*/==-10'd342+xpc10nz) || (5'd20/*MS*/==-10'd341+xpc10nz) || (5'd20/*MS*/==-10'd340+xpc10nz
              ) || (5'd20/*MS*/==-10'd338+xpc10nz) || (5'd20/*MS*/==-10'd335+xpc10nz) || (5'd20/*MS*/==-10'd334+xpc10nz) || (5'd20/*MS*/==
              -10'd330+xpc10nz) || (5'd20/*MS*/==-10'd329+xpc10nz) || (5'd20/*MS*/==-10'd327+xpc10nz) || (5'd20/*MS*/==-10'd324+xpc10nz
              ) || (5'd20/*MS*/==-10'd323+xpc10nz) || (5'd20/*MS*/==-10'd322+xpc10nz) || (5'd20/*MS*/==-10'd321+xpc10nz) || (5'd20/*MS*/==
              -10'd320+xpc10nz) || (5'd20/*MS*/==-10'd319+xpc10nz) || (5'd20/*MS*/==-10'd318+xpc10nz) || (5'd20/*MS*/==-10'd314+xpc10nz
              ) || (5'd20/*MS*/==-10'd289+xpc10nz) || (5'd20/*MS*/==-10'd287+xpc10nz) || (5'd20/*MS*/==-10'd285+xpc10nz) || (5'd20/*MS*/==
              -10'd284+xpc10nz) || (5'd20/*MS*/==-10'd259+xpc10nz) || (5'd20/*MS*/==-10'd258+xpc10nz) || (5'd20/*MS*/==-10'd257+xpc10nz
              ) || (5'd20/*MS*/==-9'd255+xpc10nz) || (5'd20/*MS*/==-9'd254+xpc10nz) || (5'd20/*MS*/==-9'd253+xpc10nz) || (5'd20/*MS*/==
              -9'd252+xpc10nz) || (5'd20/*MS*/==-9'd251+xpc10nz) || (5'd20/*MS*/==-9'd250+xpc10nz) || (5'd20/*MS*/==-9'd249+xpc10nz) || 
              (5'd20/*MS*/==-9'd248+xpc10nz) || (5'd20/*MS*/==-9'd247+xpc10nz) || (5'd20/*MS*/==-9'd246+xpc10nz) || (5'd20/*MS*/==-9'd245
              +xpc10nz) || (5'd20/*MS*/==-9'd244+xpc10nz) || (5'd20/*MS*/==-9'd242+xpc10nz) || (5'd20/*MS*/==-9'd241+xpc10nz) || (5'd20
              /*MS*/==-9'd239+xpc10nz) || (5'd20/*MS*/==-9'd238+xpc10nz) || (5'd20/*MS*/==-9'd236+xpc10nz) || (5'd20/*MS*/==-9'd171+xpc10nz
              ) || (5'd20/*MS*/==-8'd106+xpc10nz) || (5'd20/*MS*/==-8'd105+xpc10nz) || (5'd20/*MS*/==-8'd104+xpc10nz) || (5'd20/*MS*/==
              -8'd103+xpc10nz) || (5'd20/*MS*/==-8'd102+xpc10nz) || (5'd20/*MS*/==-8'd101+xpc10nz) || (5'd20/*MS*/==-8'd100+xpc10nz) || 
              (5'd20/*MS*/==-8'd99+xpc10nz) || (5'd20/*MS*/==-8'd98+xpc10nz) || (5'd20/*MS*/==-8'd97+xpc10nz) || (5'd20/*MS*/==-8'd96
              +xpc10nz) || (5'd20/*MS*/==-8'd95+xpc10nz) || (5'd20/*MS*/==-8'd94+xpc10nz) || (5'd20/*MS*/==-8'd93+xpc10nz) || (5'd20/*MS*/==
              -8'd92+xpc10nz) || (5'd20/*MS*/==-8'd91+xpc10nz) || (5'd20/*MS*/==-8'd90+xpc10nz) || (5'd20/*MS*/==-8'd89+xpc10nz) || (5'd20
              /*MS*/==-8'd88+xpc10nz) || (5'd20/*MS*/==-8'd87+xpc10nz) || (5'd20/*MS*/==-8'd86+xpc10nz) || (5'd20/*MS*/==-8'd85+xpc10nz
              ) || (5'd20/*MS*/==-8'd84+xpc10nz) || (5'd20/*MS*/==-8'd83+xpc10nz) || (5'd20/*MS*/==-8'd82+xpc10nz) || (5'd20/*MS*/==-8'd65
              +xpc10nz) || (5'd20/*MS*/==-8'd64+xpc10nz) || (5'd20/*MS*/==-7'd59+xpc10nz) || (5'd20/*MS*/==-7'd50+xpc10nz) || (5'd20/*MS*/==
              -7'd37+xpc10nz) || (5'd20/*MS*/==-6'd20+xpc10nz) || (5'd20/*MS*/==-6'd19+xpc10nz) || (5'd20/*MS*/==-6'd18+xpc10nz) || (5'd20
              /*MS*/==-6'd17+xpc10nz) || (5'd20/*MS*/==-6'd16+xpc10nz) || (5'd20/*MS*/==-5'd15+xpc10nz) || (5'd20/*MS*/==-5'd14+xpc10nz
              ) || (5'd20/*MS*/==-5'd13+xpc10nz) || (5'd20/*MS*/==-5'd12+xpc10nz) || (5'd20/*MS*/==-5'd11+xpc10nz) || (5'd20/*MS*/==-5'd10
              +xpc10nz) || (5'd20/*MS*/==-5'd9+xpc10nz) || (5'd20/*MS*/==-5'd8+xpc10nz) || (5'd20/*MS*/==-4'd7+xpc10nz) || (5'd20/*MS*/==
              -4'd6+xpc10nz) || (5'd20/*MS*/==-4'd5+xpc10nz) || (5'd20/*MS*/==-4'd4+xpc10nz) || (5'd20/*MS*/==-3'd3+xpc10nz) || (5'd20
              /*MS*/==-3'd2+xpc10nz) || (5'd20/*MS*/==-2'd1+xpc10nz) || (xpc10nz==5'd20/*US*/)) && !xpc10_clear && !xpc10_stall;

               xpc10_trk19 <= ((5'd19/*MS*/==-11'd609+xpc10nz) || (5'd19/*MS*/==-11'd599+xpc10nz) || (5'd19/*MS*/==-11'd588+xpc10nz) || 
              (5'd19/*MS*/==-11'd576+xpc10nz) || (5'd19/*MS*/==-11'd571+xpc10nz) || (5'd19/*MS*/==-11'd565+xpc10nz) || (5'd19/*MS*/==
              -11'd558+xpc10nz) || (5'd19/*MS*/==-11'd550+xpc10nz) || (5'd19/*MS*/==-11'd549+xpc10nz) || (5'd19/*MS*/==-11'd547+xpc10nz
              ) || (5'd19/*MS*/==-11'd544+xpc10nz) || (5'd19/*MS*/==-11'd540+xpc10nz) || (5'd19/*MS*/==-11'd539+xpc10nz) || (5'd19/*MS*/==
              -11'd537+xpc10nz) || (5'd19/*MS*/==-11'd534+xpc10nz) || (5'd19/*MS*/==-11'd532+xpc10nz) || (5'd19/*MS*/==-11'd528+xpc10nz
              ) || (5'd19/*MS*/==-10'd503+xpc10nz) || (5'd19/*MS*/==-10'd502+xpc10nz) || (5'd19/*MS*/==-10'd472+xpc10nz) || (5'd19/*MS*/==
              -10'd407+xpc10nz) || (5'd19/*MS*/==-10'd342+xpc10nz) || (5'd19/*MS*/==-10'd341+xpc10nz) || (5'd19/*MS*/==-10'd340+xpc10nz
              ) || (5'd19/*MS*/==-10'd338+xpc10nz) || (5'd19/*MS*/==-10'd335+xpc10nz) || (5'd19/*MS*/==-10'd334+xpc10nz) || (5'd19/*MS*/==
              -10'd330+xpc10nz) || (5'd19/*MS*/==-10'd329+xpc10nz) || (5'd19/*MS*/==-10'd327+xpc10nz) || (5'd19/*MS*/==-10'd324+xpc10nz
              ) || (5'd19/*MS*/==-10'd323+xpc10nz) || (5'd19/*MS*/==-10'd322+xpc10nz) || (5'd19/*MS*/==-10'd321+xpc10nz) || (5'd19/*MS*/==
              -10'd320+xpc10nz) || (5'd19/*MS*/==-10'd319+xpc10nz) || (5'd19/*MS*/==-10'd318+xpc10nz) || (5'd19/*MS*/==-10'd314+xpc10nz
              ) || (5'd19/*MS*/==-10'd289+xpc10nz) || (5'd19/*MS*/==-10'd287+xpc10nz) || (5'd19/*MS*/==-10'd285+xpc10nz) || (5'd19/*MS*/==
              -10'd284+xpc10nz) || (5'd19/*MS*/==-10'd259+xpc10nz) || (5'd19/*MS*/==-10'd258+xpc10nz) || (5'd19/*MS*/==-10'd257+xpc10nz
              ) || (5'd19/*MS*/==-9'd255+xpc10nz) || (5'd19/*MS*/==-9'd254+xpc10nz) || (5'd19/*MS*/==-9'd253+xpc10nz) || (5'd19/*MS*/==
              -9'd252+xpc10nz) || (5'd19/*MS*/==-9'd251+xpc10nz) || (5'd19/*MS*/==-9'd250+xpc10nz) || (5'd19/*MS*/==-9'd249+xpc10nz) || 
              (5'd19/*MS*/==-9'd248+xpc10nz) || (5'd19/*MS*/==-9'd247+xpc10nz) || (5'd19/*MS*/==-9'd246+xpc10nz) || (5'd19/*MS*/==-9'd245
              +xpc10nz) || (5'd19/*MS*/==-9'd244+xpc10nz) || (5'd19/*MS*/==-9'd242+xpc10nz) || (5'd19/*MS*/==-9'd241+xpc10nz) || (5'd19
              /*MS*/==-9'd239+xpc10nz) || (5'd19/*MS*/==-9'd238+xpc10nz) || (5'd19/*MS*/==-9'd236+xpc10nz) || (5'd19/*MS*/==-9'd171+xpc10nz
              ) || (5'd19/*MS*/==-8'd106+xpc10nz) || (5'd19/*MS*/==-8'd105+xpc10nz) || (5'd19/*MS*/==-8'd104+xpc10nz) || (5'd19/*MS*/==
              -8'd103+xpc10nz) || (5'd19/*MS*/==-8'd102+xpc10nz) || (5'd19/*MS*/==-8'd101+xpc10nz) || (5'd19/*MS*/==-8'd100+xpc10nz) || 
              (5'd19/*MS*/==-8'd99+xpc10nz) || (5'd19/*MS*/==-8'd98+xpc10nz) || (5'd19/*MS*/==-8'd97+xpc10nz) || (5'd19/*MS*/==-8'd96
              +xpc10nz) || (5'd19/*MS*/==-8'd95+xpc10nz) || (5'd19/*MS*/==-8'd94+xpc10nz) || (5'd19/*MS*/==-8'd93+xpc10nz) || (5'd19/*MS*/==
              -8'd92+xpc10nz) || (5'd19/*MS*/==-8'd91+xpc10nz) || (5'd19/*MS*/==-8'd90+xpc10nz) || (5'd19/*MS*/==-8'd89+xpc10nz) || (5'd19
              /*MS*/==-8'd88+xpc10nz) || (5'd19/*MS*/==-8'd87+xpc10nz) || (5'd19/*MS*/==-8'd86+xpc10nz) || (5'd19/*MS*/==-8'd85+xpc10nz
              ) || (5'd19/*MS*/==-8'd84+xpc10nz) || (5'd19/*MS*/==-8'd83+xpc10nz) || (5'd19/*MS*/==-8'd82+xpc10nz) || (5'd19/*MS*/==-8'd65
              +xpc10nz) || (5'd19/*MS*/==-8'd64+xpc10nz) || (5'd19/*MS*/==-7'd59+xpc10nz) || (5'd19/*MS*/==-7'd50+xpc10nz) || (5'd19/*MS*/==
              -7'd37+xpc10nz) || (5'd19/*MS*/==-6'd20+xpc10nz) || (5'd19/*MS*/==-6'd19+xpc10nz) || (5'd19/*MS*/==-6'd18+xpc10nz) || (5'd19
              /*MS*/==-6'd17+xpc10nz) || (5'd19/*MS*/==-6'd16+xpc10nz) || (5'd19/*MS*/==-5'd15+xpc10nz) || (5'd19/*MS*/==-5'd14+xpc10nz
              ) || (5'd19/*MS*/==-5'd13+xpc10nz) || (5'd19/*MS*/==-5'd12+xpc10nz) || (5'd19/*MS*/==-5'd11+xpc10nz) || (5'd19/*MS*/==-5'd10
              +xpc10nz) || (5'd19/*MS*/==-5'd9+xpc10nz) || (5'd19/*MS*/==-5'd8+xpc10nz) || (5'd19/*MS*/==-4'd7+xpc10nz) || (5'd19/*MS*/==
              -4'd6+xpc10nz) || (5'd19/*MS*/==-4'd5+xpc10nz) || (5'd19/*MS*/==-4'd4+xpc10nz) || (5'd19/*MS*/==-3'd3+xpc10nz) || (5'd19
              /*MS*/==-3'd2+xpc10nz) || (5'd19/*MS*/==-2'd1+xpc10nz) || (xpc10nz==5'd19/*US*/)) && !xpc10_clear && !xpc10_stall;

               xpc10_trk18 <= ((5'd18/*MS*/==-11'd609+xpc10nz) || (5'd18/*MS*/==-11'd599+xpc10nz) || (5'd18/*MS*/==-11'd588+xpc10nz) || 
              (5'd18/*MS*/==-11'd576+xpc10nz) || (5'd18/*MS*/==-11'd571+xpc10nz) || (5'd18/*MS*/==-11'd565+xpc10nz) || (5'd18/*MS*/==
              -11'd558+xpc10nz) || (5'd18/*MS*/==-11'd550+xpc10nz) || (5'd18/*MS*/==-11'd549+xpc10nz) || (5'd18/*MS*/==-11'd547+xpc10nz
              ) || (5'd18/*MS*/==-11'd544+xpc10nz) || (5'd18/*MS*/==-11'd540+xpc10nz) || (5'd18/*MS*/==-11'd539+xpc10nz) || (5'd18/*MS*/==
              -11'd537+xpc10nz) || (5'd18/*MS*/==-11'd534+xpc10nz) || (5'd18/*MS*/==-11'd532+xpc10nz) || (5'd18/*MS*/==-11'd528+xpc10nz
              ) || (5'd18/*MS*/==-10'd503+xpc10nz) || (5'd18/*MS*/==-10'd502+xpc10nz) || (5'd18/*MS*/==-10'd472+xpc10nz) || (5'd18/*MS*/==
              -10'd407+xpc10nz) || (5'd18/*MS*/==-10'd342+xpc10nz) || (5'd18/*MS*/==-10'd341+xpc10nz) || (5'd18/*MS*/==-10'd340+xpc10nz
              ) || (5'd18/*MS*/==-10'd338+xpc10nz) || (5'd18/*MS*/==-10'd335+xpc10nz) || (5'd18/*MS*/==-10'd334+xpc10nz) || (5'd18/*MS*/==
              -10'd330+xpc10nz) || (5'd18/*MS*/==-10'd329+xpc10nz) || (5'd18/*MS*/==-10'd327+xpc10nz) || (5'd18/*MS*/==-10'd324+xpc10nz
              ) || (5'd18/*MS*/==-10'd323+xpc10nz) || (5'd18/*MS*/==-10'd322+xpc10nz) || (5'd18/*MS*/==-10'd321+xpc10nz) || (5'd18/*MS*/==
              -10'd320+xpc10nz) || (5'd18/*MS*/==-10'd319+xpc10nz) || (5'd18/*MS*/==-10'd318+xpc10nz) || (5'd18/*MS*/==-10'd314+xpc10nz
              ) || (5'd18/*MS*/==-10'd289+xpc10nz) || (5'd18/*MS*/==-10'd287+xpc10nz) || (5'd18/*MS*/==-10'd285+xpc10nz) || (5'd18/*MS*/==
              -10'd284+xpc10nz) || (5'd18/*MS*/==-10'd259+xpc10nz) || (5'd18/*MS*/==-10'd258+xpc10nz) || (5'd18/*MS*/==-10'd257+xpc10nz
              ) || (5'd18/*MS*/==-9'd255+xpc10nz) || (5'd18/*MS*/==-9'd254+xpc10nz) || (5'd18/*MS*/==-9'd253+xpc10nz) || (5'd18/*MS*/==
              -9'd252+xpc10nz) || (5'd18/*MS*/==-9'd251+xpc10nz) || (5'd18/*MS*/==-9'd250+xpc10nz) || (5'd18/*MS*/==-9'd249+xpc10nz) || 
              (5'd18/*MS*/==-9'd248+xpc10nz) || (5'd18/*MS*/==-9'd247+xpc10nz) || (5'd18/*MS*/==-9'd246+xpc10nz) || (5'd18/*MS*/==-9'd245
              +xpc10nz) || (5'd18/*MS*/==-9'd244+xpc10nz) || (5'd18/*MS*/==-9'd242+xpc10nz) || (5'd18/*MS*/==-9'd241+xpc10nz) || (5'd18
              /*MS*/==-9'd239+xpc10nz) || (5'd18/*MS*/==-9'd238+xpc10nz) || (5'd18/*MS*/==-9'd236+xpc10nz) || (5'd18/*MS*/==-9'd171+xpc10nz
              ) || (5'd18/*MS*/==-8'd106+xpc10nz) || (5'd18/*MS*/==-8'd105+xpc10nz) || (5'd18/*MS*/==-8'd104+xpc10nz) || (5'd18/*MS*/==
              -8'd103+xpc10nz) || (5'd18/*MS*/==-8'd102+xpc10nz) || (5'd18/*MS*/==-8'd101+xpc10nz) || (5'd18/*MS*/==-8'd100+xpc10nz) || 
              (5'd18/*MS*/==-8'd99+xpc10nz) || (5'd18/*MS*/==-8'd98+xpc10nz) || (5'd18/*MS*/==-8'd97+xpc10nz) || (5'd18/*MS*/==-8'd96
              +xpc10nz) || (5'd18/*MS*/==-8'd95+xpc10nz) || (5'd18/*MS*/==-8'd94+xpc10nz) || (5'd18/*MS*/==-8'd93+xpc10nz) || (5'd18/*MS*/==
              -8'd92+xpc10nz) || (5'd18/*MS*/==-8'd91+xpc10nz) || (5'd18/*MS*/==-8'd90+xpc10nz) || (5'd18/*MS*/==-8'd89+xpc10nz) || (5'd18
              /*MS*/==-8'd88+xpc10nz) || (5'd18/*MS*/==-8'd87+xpc10nz) || (5'd18/*MS*/==-8'd86+xpc10nz) || (5'd18/*MS*/==-8'd85+xpc10nz
              ) || (5'd18/*MS*/==-8'd84+xpc10nz) || (5'd18/*MS*/==-8'd83+xpc10nz) || (5'd18/*MS*/==-8'd82+xpc10nz) || (5'd18/*MS*/==-8'd65
              +xpc10nz) || (5'd18/*MS*/==-8'd64+xpc10nz) || (5'd18/*MS*/==-7'd59+xpc10nz) || (5'd18/*MS*/==-7'd50+xpc10nz) || (5'd18/*MS*/==
              -7'd37+xpc10nz) || (5'd18/*MS*/==-6'd20+xpc10nz) || (5'd18/*MS*/==-6'd19+xpc10nz) || (5'd18/*MS*/==-6'd18+xpc10nz) || (5'd18
              /*MS*/==-6'd17+xpc10nz) || (5'd18/*MS*/==-6'd16+xpc10nz) || (5'd18/*MS*/==-5'd15+xpc10nz) || (5'd18/*MS*/==-5'd14+xpc10nz
              ) || (5'd18/*MS*/==-5'd13+xpc10nz) || (5'd18/*MS*/==-5'd12+xpc10nz) || (5'd18/*MS*/==-5'd11+xpc10nz) || (5'd18/*MS*/==-5'd10
              +xpc10nz) || (5'd18/*MS*/==-5'd9+xpc10nz) || (5'd18/*MS*/==-5'd8+xpc10nz) || (5'd18/*MS*/==-4'd7+xpc10nz) || (5'd18/*MS*/==
              -4'd6+xpc10nz) || (5'd18/*MS*/==-4'd5+xpc10nz) || (5'd18/*MS*/==-4'd4+xpc10nz) || (5'd18/*MS*/==-3'd3+xpc10nz) || (5'd18
              /*MS*/==-3'd2+xpc10nz) || (5'd18/*MS*/==-2'd1+xpc10nz) || (xpc10nz==5'd18/*US*/)) && !xpc10_clear && !xpc10_stall;

               xpc10_trk17 <= ((5'd17/*MS*/==-11'd609+xpc10nz) || (5'd17/*MS*/==-11'd599+xpc10nz) || (5'd17/*MS*/==-11'd588+xpc10nz) || 
              (5'd17/*MS*/==-11'd576+xpc10nz) || (5'd17/*MS*/==-11'd571+xpc10nz) || (5'd17/*MS*/==-11'd565+xpc10nz) || (5'd17/*MS*/==
              -11'd558+xpc10nz) || (5'd17/*MS*/==-11'd550+xpc10nz) || (5'd17/*MS*/==-11'd549+xpc10nz) || (5'd17/*MS*/==-11'd547+xpc10nz
              ) || (5'd17/*MS*/==-11'd544+xpc10nz) || (5'd17/*MS*/==-11'd540+xpc10nz) || (5'd17/*MS*/==-11'd539+xpc10nz) || (5'd17/*MS*/==
              -11'd537+xpc10nz) || (5'd17/*MS*/==-11'd534+xpc10nz) || (5'd17/*MS*/==-11'd532+xpc10nz) || (5'd17/*MS*/==-11'd528+xpc10nz
              ) || (5'd17/*MS*/==-10'd503+xpc10nz) || (5'd17/*MS*/==-10'd502+xpc10nz) || (5'd17/*MS*/==-10'd472+xpc10nz) || (5'd17/*MS*/==
              -10'd407+xpc10nz) || (5'd17/*MS*/==-10'd342+xpc10nz) || (5'd17/*MS*/==-10'd341+xpc10nz) || (5'd17/*MS*/==-10'd340+xpc10nz
              ) || (5'd17/*MS*/==-10'd338+xpc10nz) || (5'd17/*MS*/==-10'd335+xpc10nz) || (5'd17/*MS*/==-10'd334+xpc10nz) || (5'd17/*MS*/==
              -10'd330+xpc10nz) || (5'd17/*MS*/==-10'd329+xpc10nz) || (5'd17/*MS*/==-10'd327+xpc10nz) || (5'd17/*MS*/==-10'd324+xpc10nz
              ) || (5'd17/*MS*/==-10'd323+xpc10nz) || (5'd17/*MS*/==-10'd322+xpc10nz) || (5'd17/*MS*/==-10'd321+xpc10nz) || (5'd17/*MS*/==
              -10'd320+xpc10nz) || (5'd17/*MS*/==-10'd319+xpc10nz) || (5'd17/*MS*/==-10'd318+xpc10nz) || (5'd17/*MS*/==-10'd314+xpc10nz
              ) || (5'd17/*MS*/==-10'd289+xpc10nz) || (5'd17/*MS*/==-10'd287+xpc10nz) || (5'd17/*MS*/==-10'd285+xpc10nz) || (5'd17/*MS*/==
              -10'd284+xpc10nz) || (5'd17/*MS*/==-10'd259+xpc10nz) || (5'd17/*MS*/==-10'd258+xpc10nz) || (5'd17/*MS*/==-10'd257+xpc10nz
              ) || (5'd17/*MS*/==-9'd255+xpc10nz) || (5'd17/*MS*/==-9'd254+xpc10nz) || (5'd17/*MS*/==-9'd253+xpc10nz) || (5'd17/*MS*/==
              -9'd252+xpc10nz) || (5'd17/*MS*/==-9'd251+xpc10nz) || (5'd17/*MS*/==-9'd250+xpc10nz) || (5'd17/*MS*/==-9'd249+xpc10nz) || 
              (5'd17/*MS*/==-9'd248+xpc10nz) || (5'd17/*MS*/==-9'd247+xpc10nz) || (5'd17/*MS*/==-9'd246+xpc10nz) || (5'd17/*MS*/==-9'd245
              +xpc10nz) || (5'd17/*MS*/==-9'd244+xpc10nz) || (5'd17/*MS*/==-9'd242+xpc10nz) || (5'd17/*MS*/==-9'd241+xpc10nz) || (5'd17
              /*MS*/==-9'd239+xpc10nz) || (5'd17/*MS*/==-9'd238+xpc10nz) || (5'd17/*MS*/==-9'd236+xpc10nz) || (5'd17/*MS*/==-9'd171+xpc10nz
              ) || (5'd17/*MS*/==-8'd106+xpc10nz) || (5'd17/*MS*/==-8'd105+xpc10nz) || (5'd17/*MS*/==-8'd104+xpc10nz) || (5'd17/*MS*/==
              -8'd103+xpc10nz) || (5'd17/*MS*/==-8'd102+xpc10nz) || (5'd17/*MS*/==-8'd101+xpc10nz) || (5'd17/*MS*/==-8'd100+xpc10nz) || 
              (5'd17/*MS*/==-8'd99+xpc10nz) || (5'd17/*MS*/==-8'd98+xpc10nz) || (5'd17/*MS*/==-8'd97+xpc10nz) || (5'd17/*MS*/==-8'd96
              +xpc10nz) || (5'd17/*MS*/==-8'd95+xpc10nz) || (5'd17/*MS*/==-8'd94+xpc10nz) || (5'd17/*MS*/==-8'd93+xpc10nz) || (5'd17/*MS*/==
              -8'd92+xpc10nz) || (5'd17/*MS*/==-8'd91+xpc10nz) || (5'd17/*MS*/==-8'd90+xpc10nz) || (5'd17/*MS*/==-8'd89+xpc10nz) || (5'd17
              /*MS*/==-8'd88+xpc10nz) || (5'd17/*MS*/==-8'd87+xpc10nz) || (5'd17/*MS*/==-8'd86+xpc10nz) || (5'd17/*MS*/==-8'd85+xpc10nz
              ) || (5'd17/*MS*/==-8'd84+xpc10nz) || (5'd17/*MS*/==-8'd83+xpc10nz) || (5'd17/*MS*/==-8'd82+xpc10nz) || (5'd17/*MS*/==-8'd65
              +xpc10nz) || (5'd17/*MS*/==-8'd64+xpc10nz) || (5'd17/*MS*/==-7'd59+xpc10nz) || (5'd17/*MS*/==-7'd50+xpc10nz) || (5'd17/*MS*/==
              -7'd37+xpc10nz) || (5'd17/*MS*/==-6'd20+xpc10nz) || (5'd17/*MS*/==-6'd19+xpc10nz) || (5'd17/*MS*/==-6'd18+xpc10nz) || (5'd17
              /*MS*/==-6'd17+xpc10nz) || (5'd17/*MS*/==-6'd16+xpc10nz) || (5'd17/*MS*/==-5'd15+xpc10nz) || (5'd17/*MS*/==-5'd14+xpc10nz
              ) || (5'd17/*MS*/==-5'd13+xpc10nz) || (5'd17/*MS*/==-5'd12+xpc10nz) || (5'd17/*MS*/==-5'd11+xpc10nz) || (5'd17/*MS*/==-5'd10
              +xpc10nz) || (5'd17/*MS*/==-5'd9+xpc10nz) || (5'd17/*MS*/==-5'd8+xpc10nz) || (5'd17/*MS*/==-4'd7+xpc10nz) || (5'd17/*MS*/==
              -4'd6+xpc10nz) || (5'd17/*MS*/==-4'd5+xpc10nz) || (5'd17/*MS*/==-4'd4+xpc10nz) || (5'd17/*MS*/==-3'd3+xpc10nz) || (5'd17
              /*MS*/==-3'd2+xpc10nz) || (5'd17/*MS*/==-2'd1+xpc10nz) || (xpc10nz==5'd17/*US*/)) && !xpc10_clear && !xpc10_stall;

               xpc10_trk16 <= ((5'd16/*MS*/==-11'd609+xpc10nz) || (5'd16/*MS*/==-11'd599+xpc10nz) || (5'd16/*MS*/==-11'd588+xpc10nz) || 
              (5'd16/*MS*/==-11'd576+xpc10nz) || (5'd16/*MS*/==-11'd571+xpc10nz) || (5'd16/*MS*/==-11'd565+xpc10nz) || (5'd16/*MS*/==
              -11'd558+xpc10nz) || (5'd16/*MS*/==-11'd550+xpc10nz) || (5'd16/*MS*/==-11'd549+xpc10nz) || (5'd16/*MS*/==-11'd547+xpc10nz
              ) || (5'd16/*MS*/==-11'd544+xpc10nz) || (5'd16/*MS*/==-11'd540+xpc10nz) || (5'd16/*MS*/==-11'd539+xpc10nz) || (5'd16/*MS*/==
              -11'd537+xpc10nz) || (5'd16/*MS*/==-11'd534+xpc10nz) || (5'd16/*MS*/==-11'd532+xpc10nz) || (5'd16/*MS*/==-11'd528+xpc10nz
              ) || (5'd16/*MS*/==-10'd503+xpc10nz) || (5'd16/*MS*/==-10'd502+xpc10nz) || (5'd16/*MS*/==-10'd472+xpc10nz) || (5'd16/*MS*/==
              -10'd407+xpc10nz) || (5'd16/*MS*/==-10'd342+xpc10nz) || (5'd16/*MS*/==-10'd341+xpc10nz) || (5'd16/*MS*/==-10'd340+xpc10nz
              ) || (5'd16/*MS*/==-10'd338+xpc10nz) || (5'd16/*MS*/==-10'd335+xpc10nz) || (5'd16/*MS*/==-10'd334+xpc10nz) || (5'd16/*MS*/==
              -10'd330+xpc10nz) || (5'd16/*MS*/==-10'd329+xpc10nz) || (5'd16/*MS*/==-10'd327+xpc10nz) || (5'd16/*MS*/==-10'd324+xpc10nz
              ) || (5'd16/*MS*/==-10'd323+xpc10nz) || (5'd16/*MS*/==-10'd322+xpc10nz) || (5'd16/*MS*/==-10'd321+xpc10nz) || (5'd16/*MS*/==
              -10'd320+xpc10nz) || (5'd16/*MS*/==-10'd319+xpc10nz) || (5'd16/*MS*/==-10'd318+xpc10nz) || (5'd16/*MS*/==-10'd314+xpc10nz
              ) || (5'd16/*MS*/==-10'd289+xpc10nz) || (5'd16/*MS*/==-10'd287+xpc10nz) || (5'd16/*MS*/==-10'd285+xpc10nz) || (5'd16/*MS*/==
              -10'd284+xpc10nz) || (5'd16/*MS*/==-10'd259+xpc10nz) || (5'd16/*MS*/==-10'd258+xpc10nz) || (5'd16/*MS*/==-10'd257+xpc10nz
              ) || (5'd16/*MS*/==-9'd255+xpc10nz) || (5'd16/*MS*/==-9'd254+xpc10nz) || (5'd16/*MS*/==-9'd253+xpc10nz) || (5'd16/*MS*/==
              -9'd252+xpc10nz) || (5'd16/*MS*/==-9'd251+xpc10nz) || (5'd16/*MS*/==-9'd250+xpc10nz) || (5'd16/*MS*/==-9'd249+xpc10nz) || 
              (5'd16/*MS*/==-9'd248+xpc10nz) || (5'd16/*MS*/==-9'd247+xpc10nz) || (5'd16/*MS*/==-9'd246+xpc10nz) || (5'd16/*MS*/==-9'd245
              +xpc10nz) || (5'd16/*MS*/==-9'd244+xpc10nz) || (5'd16/*MS*/==-9'd242+xpc10nz) || (5'd16/*MS*/==-9'd241+xpc10nz) || (5'd16
              /*MS*/==-9'd239+xpc10nz) || (5'd16/*MS*/==-9'd238+xpc10nz) || (5'd16/*MS*/==-9'd236+xpc10nz) || (5'd16/*MS*/==-9'd171+xpc10nz
              ) || (5'd16/*MS*/==-8'd106+xpc10nz) || (5'd16/*MS*/==-8'd105+xpc10nz) || (5'd16/*MS*/==-8'd104+xpc10nz) || (5'd16/*MS*/==
              -8'd103+xpc10nz) || (5'd16/*MS*/==-8'd102+xpc10nz) || (5'd16/*MS*/==-8'd101+xpc10nz) || (5'd16/*MS*/==-8'd100+xpc10nz) || 
              (5'd16/*MS*/==-8'd99+xpc10nz) || (5'd16/*MS*/==-8'd98+xpc10nz) || (5'd16/*MS*/==-8'd97+xpc10nz) || (5'd16/*MS*/==-8'd96
              +xpc10nz) || (5'd16/*MS*/==-8'd95+xpc10nz) || (5'd16/*MS*/==-8'd94+xpc10nz) || (5'd16/*MS*/==-8'd93+xpc10nz) || (5'd16/*MS*/==
              -8'd92+xpc10nz) || (5'd16/*MS*/==-8'd91+xpc10nz) || (5'd16/*MS*/==-8'd90+xpc10nz) || (5'd16/*MS*/==-8'd89+xpc10nz) || (5'd16
              /*MS*/==-8'd88+xpc10nz) || (5'd16/*MS*/==-8'd87+xpc10nz) || (5'd16/*MS*/==-8'd86+xpc10nz) || (5'd16/*MS*/==-8'd85+xpc10nz
              ) || (5'd16/*MS*/==-8'd84+xpc10nz) || (5'd16/*MS*/==-8'd83+xpc10nz) || (5'd16/*MS*/==-8'd82+xpc10nz) || (5'd16/*MS*/==-8'd65
              +xpc10nz) || (5'd16/*MS*/==-8'd64+xpc10nz) || (5'd16/*MS*/==-7'd59+xpc10nz) || (5'd16/*MS*/==-7'd50+xpc10nz) || (5'd16/*MS*/==
              -7'd37+xpc10nz) || (5'd16/*MS*/==-6'd20+xpc10nz) || (5'd16/*MS*/==-6'd19+xpc10nz) || (5'd16/*MS*/==-6'd18+xpc10nz) || (5'd16
              /*MS*/==-6'd17+xpc10nz) || (5'd16/*MS*/==-6'd16+xpc10nz) || (5'd16/*MS*/==-5'd15+xpc10nz) || (5'd16/*MS*/==-5'd14+xpc10nz
              ) || (5'd16/*MS*/==-5'd13+xpc10nz) || (5'd16/*MS*/==-5'd12+xpc10nz) || (5'd16/*MS*/==-5'd11+xpc10nz) || (5'd16/*MS*/==-5'd10
              +xpc10nz) || (5'd16/*MS*/==-5'd9+xpc10nz) || (5'd16/*MS*/==-5'd8+xpc10nz) || (5'd16/*MS*/==-4'd7+xpc10nz) || (5'd16/*MS*/==
              -4'd6+xpc10nz) || (5'd16/*MS*/==-4'd5+xpc10nz) || (5'd16/*MS*/==-4'd4+xpc10nz) || (5'd16/*MS*/==-3'd3+xpc10nz) || (5'd16
              /*MS*/==-3'd2+xpc10nz) || (5'd16/*MS*/==-2'd1+xpc10nz) || (xpc10nz==5'd16/*US*/)) && !xpc10_clear && !xpc10_stall;

               xpc10_trk15 <= ((4'd15/*MS*/==-11'd609+xpc10nz) || (4'd15/*MS*/==-11'd599+xpc10nz) || (4'd15/*MS*/==-11'd588+xpc10nz) || 
              (4'd15/*MS*/==-11'd576+xpc10nz) || (4'd15/*MS*/==-11'd571+xpc10nz) || (4'd15/*MS*/==-11'd565+xpc10nz) || (4'd15/*MS*/==
              -11'd558+xpc10nz) || (4'd15/*MS*/==-11'd550+xpc10nz) || (4'd15/*MS*/==-11'd549+xpc10nz) || (4'd15/*MS*/==-11'd547+xpc10nz
              ) || (4'd15/*MS*/==-11'd544+xpc10nz) || (4'd15/*MS*/==-11'd540+xpc10nz) || (4'd15/*MS*/==-11'd539+xpc10nz) || (4'd15/*MS*/==
              -11'd537+xpc10nz) || (4'd15/*MS*/==-11'd534+xpc10nz) || (4'd15/*MS*/==-11'd532+xpc10nz) || (4'd15/*MS*/==-11'd528+xpc10nz
              ) || (4'd15/*MS*/==-10'd503+xpc10nz) || (4'd15/*MS*/==-10'd502+xpc10nz) || (4'd15/*MS*/==-10'd472+xpc10nz) || (4'd15/*MS*/==
              -10'd407+xpc10nz) || (4'd15/*MS*/==-10'd342+xpc10nz) || (4'd15/*MS*/==-10'd341+xpc10nz) || (4'd15/*MS*/==-10'd340+xpc10nz
              ) || (4'd15/*MS*/==-10'd338+xpc10nz) || (4'd15/*MS*/==-10'd335+xpc10nz) || (4'd15/*MS*/==-10'd334+xpc10nz) || (4'd15/*MS*/==
              -10'd330+xpc10nz) || (4'd15/*MS*/==-10'd329+xpc10nz) || (4'd15/*MS*/==-10'd327+xpc10nz) || (4'd15/*MS*/==-10'd324+xpc10nz
              ) || (4'd15/*MS*/==-10'd323+xpc10nz) || (4'd15/*MS*/==-10'd322+xpc10nz) || (4'd15/*MS*/==-10'd321+xpc10nz) || (4'd15/*MS*/==
              -10'd320+xpc10nz) || (4'd15/*MS*/==-10'd319+xpc10nz) || (4'd15/*MS*/==-10'd318+xpc10nz) || (4'd15/*MS*/==-10'd314+xpc10nz
              ) || (4'd15/*MS*/==-10'd289+xpc10nz) || (4'd15/*MS*/==-10'd287+xpc10nz) || (4'd15/*MS*/==-10'd285+xpc10nz) || (4'd15/*MS*/==
              -10'd284+xpc10nz) || (4'd15/*MS*/==-10'd259+xpc10nz) || (4'd15/*MS*/==-10'd258+xpc10nz) || (4'd15/*MS*/==-10'd257+xpc10nz
              ) || (4'd15/*MS*/==-9'd255+xpc10nz) || (4'd15/*MS*/==-9'd254+xpc10nz) || (4'd15/*MS*/==-9'd253+xpc10nz) || (4'd15/*MS*/==
              -9'd252+xpc10nz) || (4'd15/*MS*/==-9'd251+xpc10nz) || (4'd15/*MS*/==-9'd250+xpc10nz) || (4'd15/*MS*/==-9'd249+xpc10nz) || 
              (4'd15/*MS*/==-9'd248+xpc10nz) || (4'd15/*MS*/==-9'd247+xpc10nz) || (4'd15/*MS*/==-9'd246+xpc10nz) || (4'd15/*MS*/==-9'd245
              +xpc10nz) || (4'd15/*MS*/==-9'd244+xpc10nz) || (4'd15/*MS*/==-9'd242+xpc10nz) || (4'd15/*MS*/==-9'd241+xpc10nz) || (4'd15
              /*MS*/==-9'd239+xpc10nz) || (4'd15/*MS*/==-9'd238+xpc10nz) || (4'd15/*MS*/==-9'd236+xpc10nz) || (4'd15/*MS*/==-9'd171+xpc10nz
              ) || (4'd15/*MS*/==-8'd106+xpc10nz) || (4'd15/*MS*/==-8'd105+xpc10nz) || (4'd15/*MS*/==-8'd104+xpc10nz) || (4'd15/*MS*/==
              -8'd103+xpc10nz) || (4'd15/*MS*/==-8'd102+xpc10nz) || (4'd15/*MS*/==-8'd101+xpc10nz) || (4'd15/*MS*/==-8'd100+xpc10nz) || 
              (4'd15/*MS*/==-8'd99+xpc10nz) || (4'd15/*MS*/==-8'd98+xpc10nz) || (4'd15/*MS*/==-8'd97+xpc10nz) || (4'd15/*MS*/==-8'd96
              +xpc10nz) || (4'd15/*MS*/==-8'd95+xpc10nz) || (4'd15/*MS*/==-8'd94+xpc10nz) || (4'd15/*MS*/==-8'd93+xpc10nz) || (4'd15/*MS*/==
              -8'd92+xpc10nz) || (4'd15/*MS*/==-8'd91+xpc10nz) || (4'd15/*MS*/==-8'd90+xpc10nz) || (4'd15/*MS*/==-8'd89+xpc10nz) || (4'd15
              /*MS*/==-8'd88+xpc10nz) || (4'd15/*MS*/==-8'd87+xpc10nz) || (4'd15/*MS*/==-8'd86+xpc10nz) || (4'd15/*MS*/==-8'd85+xpc10nz
              ) || (4'd15/*MS*/==-8'd84+xpc10nz) || (4'd15/*MS*/==-8'd83+xpc10nz) || (4'd15/*MS*/==-8'd82+xpc10nz) || (4'd15/*MS*/==-8'd65
              +xpc10nz) || (4'd15/*MS*/==-8'd64+xpc10nz) || (4'd15/*MS*/==-7'd59+xpc10nz) || (4'd15/*MS*/==-7'd50+xpc10nz) || (4'd15/*MS*/==
              -7'd37+xpc10nz) || (4'd15/*MS*/==-6'd20+xpc10nz) || (4'd15/*MS*/==-6'd19+xpc10nz) || (4'd15/*MS*/==-6'd18+xpc10nz) || (4'd15
              /*MS*/==-6'd17+xpc10nz) || (4'd15/*MS*/==-6'd16+xpc10nz) || (4'd15/*MS*/==-5'd15+xpc10nz) || (4'd15/*MS*/==-5'd14+xpc10nz
              ) || (4'd15/*MS*/==-5'd13+xpc10nz) || (4'd15/*MS*/==-5'd12+xpc10nz) || (4'd15/*MS*/==-5'd11+xpc10nz) || (4'd15/*MS*/==-5'd10
              +xpc10nz) || (4'd15/*MS*/==-5'd9+xpc10nz) || (4'd15/*MS*/==-5'd8+xpc10nz) || (4'd15/*MS*/==-4'd7+xpc10nz) || (4'd15/*MS*/==
              -4'd6+xpc10nz) || (4'd15/*MS*/==-4'd5+xpc10nz) || (4'd15/*MS*/==-4'd4+xpc10nz) || (4'd15/*MS*/==-3'd3+xpc10nz) || (4'd15
              /*MS*/==-3'd2+xpc10nz) || (4'd15/*MS*/==-2'd1+xpc10nz) || (xpc10nz==4'd15/*US*/)) && !xpc10_clear && !xpc10_stall;

               xpc10_trk14 <= ((4'd14/*MS*/==-11'd609+xpc10nz) || (4'd14/*MS*/==-11'd599+xpc10nz) || (4'd14/*MS*/==-11'd588+xpc10nz) || 
              (4'd14/*MS*/==-11'd576+xpc10nz) || (4'd14/*MS*/==-11'd571+xpc10nz) || (4'd14/*MS*/==-11'd565+xpc10nz) || (4'd14/*MS*/==
              -11'd558+xpc10nz) || (4'd14/*MS*/==-11'd550+xpc10nz) || (4'd14/*MS*/==-11'd549+xpc10nz) || (4'd14/*MS*/==-11'd547+xpc10nz
              ) || (4'd14/*MS*/==-11'd544+xpc10nz) || (4'd14/*MS*/==-11'd540+xpc10nz) || (4'd14/*MS*/==-11'd539+xpc10nz) || (4'd14/*MS*/==
              -11'd537+xpc10nz) || (4'd14/*MS*/==-11'd534+xpc10nz) || (4'd14/*MS*/==-11'd532+xpc10nz) || (4'd14/*MS*/==-11'd528+xpc10nz
              ) || (4'd14/*MS*/==-10'd503+xpc10nz) || (4'd14/*MS*/==-10'd502+xpc10nz) || (4'd14/*MS*/==-10'd472+xpc10nz) || (4'd14/*MS*/==
              -10'd407+xpc10nz) || (4'd14/*MS*/==-10'd342+xpc10nz) || (4'd14/*MS*/==-10'd341+xpc10nz) || (4'd14/*MS*/==-10'd340+xpc10nz
              ) || (4'd14/*MS*/==-10'd338+xpc10nz) || (4'd14/*MS*/==-10'd335+xpc10nz) || (4'd14/*MS*/==-10'd334+xpc10nz) || (4'd14/*MS*/==
              -10'd330+xpc10nz) || (4'd14/*MS*/==-10'd329+xpc10nz) || (4'd14/*MS*/==-10'd327+xpc10nz) || (4'd14/*MS*/==-10'd324+xpc10nz
              ) || (4'd14/*MS*/==-10'd323+xpc10nz) || (4'd14/*MS*/==-10'd322+xpc10nz) || (4'd14/*MS*/==-10'd321+xpc10nz) || (4'd14/*MS*/==
              -10'd320+xpc10nz) || (4'd14/*MS*/==-10'd319+xpc10nz) || (4'd14/*MS*/==-10'd318+xpc10nz) || (4'd14/*MS*/==-10'd314+xpc10nz
              ) || (4'd14/*MS*/==-10'd289+xpc10nz) || (4'd14/*MS*/==-10'd287+xpc10nz) || (4'd14/*MS*/==-10'd285+xpc10nz) || (4'd14/*MS*/==
              -10'd284+xpc10nz) || (4'd14/*MS*/==-10'd259+xpc10nz) || (4'd14/*MS*/==-10'd258+xpc10nz) || (4'd14/*MS*/==-10'd257+xpc10nz
              ) || (4'd14/*MS*/==-9'd255+xpc10nz) || (4'd14/*MS*/==-9'd254+xpc10nz) || (4'd14/*MS*/==-9'd253+xpc10nz) || (4'd14/*MS*/==
              -9'd252+xpc10nz) || (4'd14/*MS*/==-9'd251+xpc10nz) || (4'd14/*MS*/==-9'd250+xpc10nz) || (4'd14/*MS*/==-9'd249+xpc10nz) || 
              (4'd14/*MS*/==-9'd248+xpc10nz) || (4'd14/*MS*/==-9'd247+xpc10nz) || (4'd14/*MS*/==-9'd246+xpc10nz) || (4'd14/*MS*/==-9'd245
              +xpc10nz) || (4'd14/*MS*/==-9'd244+xpc10nz) || (4'd14/*MS*/==-9'd242+xpc10nz) || (4'd14/*MS*/==-9'd241+xpc10nz) || (4'd14
              /*MS*/==-9'd239+xpc10nz) || (4'd14/*MS*/==-9'd238+xpc10nz) || (4'd14/*MS*/==-9'd236+xpc10nz) || (4'd14/*MS*/==-9'd171+xpc10nz
              ) || (4'd14/*MS*/==-8'd106+xpc10nz) || (4'd14/*MS*/==-8'd105+xpc10nz) || (4'd14/*MS*/==-8'd104+xpc10nz) || (4'd14/*MS*/==
              -8'd103+xpc10nz) || (4'd14/*MS*/==-8'd102+xpc10nz) || (4'd14/*MS*/==-8'd101+xpc10nz) || (4'd14/*MS*/==-8'd100+xpc10nz) || 
              (4'd14/*MS*/==-8'd99+xpc10nz) || (4'd14/*MS*/==-8'd98+xpc10nz) || (4'd14/*MS*/==-8'd97+xpc10nz) || (4'd14/*MS*/==-8'd96
              +xpc10nz) || (4'd14/*MS*/==-8'd95+xpc10nz) || (4'd14/*MS*/==-8'd94+xpc10nz) || (4'd14/*MS*/==-8'd93+xpc10nz) || (4'd14/*MS*/==
              -8'd92+xpc10nz) || (4'd14/*MS*/==-8'd91+xpc10nz) || (4'd14/*MS*/==-8'd90+xpc10nz) || (4'd14/*MS*/==-8'd89+xpc10nz) || (4'd14
              /*MS*/==-8'd88+xpc10nz) || (4'd14/*MS*/==-8'd87+xpc10nz) || (4'd14/*MS*/==-8'd86+xpc10nz) || (4'd14/*MS*/==-8'd85+xpc10nz
              ) || (4'd14/*MS*/==-8'd84+xpc10nz) || (4'd14/*MS*/==-8'd83+xpc10nz) || (4'd14/*MS*/==-8'd82+xpc10nz) || (4'd14/*MS*/==-8'd65
              +xpc10nz) || (4'd14/*MS*/==-8'd64+xpc10nz) || (4'd14/*MS*/==-7'd59+xpc10nz) || (4'd14/*MS*/==-7'd50+xpc10nz) || (4'd14/*MS*/==
              -7'd37+xpc10nz) || (4'd14/*MS*/==-6'd20+xpc10nz) || (4'd14/*MS*/==-6'd19+xpc10nz) || (4'd14/*MS*/==-6'd18+xpc10nz) || (4'd14
              /*MS*/==-6'd17+xpc10nz) || (4'd14/*MS*/==-6'd16+xpc10nz) || (4'd14/*MS*/==-5'd15+xpc10nz) || (4'd14/*MS*/==-5'd14+xpc10nz
              ) || (4'd14/*MS*/==-5'd13+xpc10nz) || (4'd14/*MS*/==-5'd12+xpc10nz) || (4'd14/*MS*/==-5'd11+xpc10nz) || (4'd14/*MS*/==-5'd10
              +xpc10nz) || (4'd14/*MS*/==-5'd9+xpc10nz) || (4'd14/*MS*/==-5'd8+xpc10nz) || (4'd14/*MS*/==-4'd7+xpc10nz) || (4'd14/*MS*/==
              -4'd6+xpc10nz) || (4'd14/*MS*/==-4'd5+xpc10nz) || (4'd14/*MS*/==-4'd4+xpc10nz) || (4'd14/*MS*/==-3'd3+xpc10nz) || (4'd14
              /*MS*/==-3'd2+xpc10nz) || (4'd14/*MS*/==-2'd1+xpc10nz) || (xpc10nz==4'd14/*US*/)) && !xpc10_clear && !xpc10_stall;

               xpc10_trk13 <= ((4'd13/*MS*/==-11'd609+xpc10nz) || (4'd13/*MS*/==-11'd599+xpc10nz) || (4'd13/*MS*/==-11'd588+xpc10nz) || 
              (4'd13/*MS*/==-11'd576+xpc10nz) || (4'd13/*MS*/==-11'd571+xpc10nz) || (4'd13/*MS*/==-11'd565+xpc10nz) || (4'd13/*MS*/==
              -11'd558+xpc10nz) || (4'd13/*MS*/==-11'd550+xpc10nz) || (4'd13/*MS*/==-11'd549+xpc10nz) || (4'd13/*MS*/==-11'd547+xpc10nz
              ) || (4'd13/*MS*/==-11'd544+xpc10nz) || (4'd13/*MS*/==-11'd540+xpc10nz) || (4'd13/*MS*/==-11'd539+xpc10nz) || (4'd13/*MS*/==
              -11'd537+xpc10nz) || (4'd13/*MS*/==-11'd534+xpc10nz) || (4'd13/*MS*/==-11'd532+xpc10nz) || (4'd13/*MS*/==-11'd528+xpc10nz
              ) || (4'd13/*MS*/==-10'd503+xpc10nz) || (4'd13/*MS*/==-10'd502+xpc10nz) || (4'd13/*MS*/==-10'd472+xpc10nz) || (4'd13/*MS*/==
              -10'd407+xpc10nz) || (4'd13/*MS*/==-10'd342+xpc10nz) || (4'd13/*MS*/==-10'd341+xpc10nz) || (4'd13/*MS*/==-10'd340+xpc10nz
              ) || (4'd13/*MS*/==-10'd338+xpc10nz) || (4'd13/*MS*/==-10'd335+xpc10nz) || (4'd13/*MS*/==-10'd334+xpc10nz) || (4'd13/*MS*/==
              -10'd330+xpc10nz) || (4'd13/*MS*/==-10'd329+xpc10nz) || (4'd13/*MS*/==-10'd327+xpc10nz) || (4'd13/*MS*/==-10'd324+xpc10nz
              ) || (4'd13/*MS*/==-10'd323+xpc10nz) || (4'd13/*MS*/==-10'd322+xpc10nz) || (4'd13/*MS*/==-10'd321+xpc10nz) || (4'd13/*MS*/==
              -10'd320+xpc10nz) || (4'd13/*MS*/==-10'd319+xpc10nz) || (4'd13/*MS*/==-10'd318+xpc10nz) || (4'd13/*MS*/==-10'd314+xpc10nz
              ) || (4'd13/*MS*/==-10'd289+xpc10nz) || (4'd13/*MS*/==-10'd287+xpc10nz) || (4'd13/*MS*/==-10'd285+xpc10nz) || (4'd13/*MS*/==
              -10'd284+xpc10nz) || (4'd13/*MS*/==-10'd259+xpc10nz) || (4'd13/*MS*/==-10'd258+xpc10nz) || (4'd13/*MS*/==-10'd257+xpc10nz
              ) || (4'd13/*MS*/==-9'd255+xpc10nz) || (4'd13/*MS*/==-9'd254+xpc10nz) || (4'd13/*MS*/==-9'd253+xpc10nz) || (4'd13/*MS*/==
              -9'd252+xpc10nz) || (4'd13/*MS*/==-9'd251+xpc10nz) || (4'd13/*MS*/==-9'd250+xpc10nz) || (4'd13/*MS*/==-9'd249+xpc10nz) || 
              (4'd13/*MS*/==-9'd248+xpc10nz) || (4'd13/*MS*/==-9'd247+xpc10nz) || (4'd13/*MS*/==-9'd246+xpc10nz) || (4'd13/*MS*/==-9'd245
              +xpc10nz) || (4'd13/*MS*/==-9'd244+xpc10nz) || (4'd13/*MS*/==-9'd242+xpc10nz) || (4'd13/*MS*/==-9'd241+xpc10nz) || (4'd13
              /*MS*/==-9'd239+xpc10nz) || (4'd13/*MS*/==-9'd238+xpc10nz) || (4'd13/*MS*/==-9'd236+xpc10nz) || (4'd13/*MS*/==-9'd171+xpc10nz
              ) || (4'd13/*MS*/==-8'd106+xpc10nz) || (4'd13/*MS*/==-8'd105+xpc10nz) || (4'd13/*MS*/==-8'd104+xpc10nz) || (4'd13/*MS*/==
              -8'd103+xpc10nz) || (4'd13/*MS*/==-8'd102+xpc10nz) || (4'd13/*MS*/==-8'd101+xpc10nz) || (4'd13/*MS*/==-8'd100+xpc10nz) || 
              (4'd13/*MS*/==-8'd99+xpc10nz) || (4'd13/*MS*/==-8'd98+xpc10nz) || (4'd13/*MS*/==-8'd97+xpc10nz) || (4'd13/*MS*/==-8'd96
              +xpc10nz) || (4'd13/*MS*/==-8'd95+xpc10nz) || (4'd13/*MS*/==-8'd94+xpc10nz) || (4'd13/*MS*/==-8'd93+xpc10nz) || (4'd13/*MS*/==
              -8'd92+xpc10nz) || (4'd13/*MS*/==-8'd91+xpc10nz) || (4'd13/*MS*/==-8'd90+xpc10nz) || (4'd13/*MS*/==-8'd89+xpc10nz) || (4'd13
              /*MS*/==-8'd88+xpc10nz) || (4'd13/*MS*/==-8'd87+xpc10nz) || (4'd13/*MS*/==-8'd86+xpc10nz) || (4'd13/*MS*/==-8'd85+xpc10nz
              ) || (4'd13/*MS*/==-8'd84+xpc10nz) || (4'd13/*MS*/==-8'd83+xpc10nz) || (4'd13/*MS*/==-8'd82+xpc10nz) || (4'd13/*MS*/==-8'd65
              +xpc10nz) || (4'd13/*MS*/==-8'd64+xpc10nz) || (4'd13/*MS*/==-7'd59+xpc10nz) || (4'd13/*MS*/==-7'd50+xpc10nz) || (4'd13/*MS*/==
              -7'd37+xpc10nz) || (4'd13/*MS*/==-6'd20+xpc10nz) || (4'd13/*MS*/==-6'd19+xpc10nz) || (4'd13/*MS*/==-6'd18+xpc10nz) || (4'd13
              /*MS*/==-6'd17+xpc10nz) || (4'd13/*MS*/==-6'd16+xpc10nz) || (4'd13/*MS*/==-5'd15+xpc10nz) || (4'd13/*MS*/==-5'd14+xpc10nz
              ) || (4'd13/*MS*/==-5'd13+xpc10nz) || (4'd13/*MS*/==-5'd12+xpc10nz) || (4'd13/*MS*/==-5'd11+xpc10nz) || (4'd13/*MS*/==-5'd10
              +xpc10nz) || (4'd13/*MS*/==-5'd9+xpc10nz) || (4'd13/*MS*/==-5'd8+xpc10nz) || (4'd13/*MS*/==-4'd7+xpc10nz) || (4'd13/*MS*/==
              -4'd6+xpc10nz) || (4'd13/*MS*/==-4'd5+xpc10nz) || (4'd13/*MS*/==-4'd4+xpc10nz) || (4'd13/*MS*/==-3'd3+xpc10nz) || (4'd13
              /*MS*/==-3'd2+xpc10nz) || (4'd13/*MS*/==-2'd1+xpc10nz) || (xpc10nz==4'd13/*US*/)) && !xpc10_clear && !xpc10_stall;

               xpc10_trk12 <= ((4'd12/*MS*/==-11'd609+xpc10nz) || (4'd12/*MS*/==-11'd599+xpc10nz) || (4'd12/*MS*/==-11'd588+xpc10nz) || 
              (4'd12/*MS*/==-11'd576+xpc10nz) || (4'd12/*MS*/==-11'd571+xpc10nz) || (4'd12/*MS*/==-11'd565+xpc10nz) || (4'd12/*MS*/==
              -11'd558+xpc10nz) || (4'd12/*MS*/==-11'd550+xpc10nz) || (4'd12/*MS*/==-11'd549+xpc10nz) || (4'd12/*MS*/==-11'd547+xpc10nz
              ) || (4'd12/*MS*/==-11'd544+xpc10nz) || (4'd12/*MS*/==-11'd540+xpc10nz) || (4'd12/*MS*/==-11'd539+xpc10nz) || (4'd12/*MS*/==
              -11'd537+xpc10nz) || (4'd12/*MS*/==-11'd534+xpc10nz) || (4'd12/*MS*/==-11'd532+xpc10nz) || (4'd12/*MS*/==-11'd528+xpc10nz
              ) || (4'd12/*MS*/==-10'd503+xpc10nz) || (4'd12/*MS*/==-10'd502+xpc10nz) || (4'd12/*MS*/==-10'd472+xpc10nz) || (4'd12/*MS*/==
              -10'd407+xpc10nz) || (4'd12/*MS*/==-10'd342+xpc10nz) || (4'd12/*MS*/==-10'd341+xpc10nz) || (4'd12/*MS*/==-10'd340+xpc10nz
              ) || (4'd12/*MS*/==-10'd338+xpc10nz) || (4'd12/*MS*/==-10'd335+xpc10nz) || (4'd12/*MS*/==-10'd334+xpc10nz) || (4'd12/*MS*/==
              -10'd330+xpc10nz) || (4'd12/*MS*/==-10'd329+xpc10nz) || (4'd12/*MS*/==-10'd327+xpc10nz) || (4'd12/*MS*/==-10'd324+xpc10nz
              ) || (4'd12/*MS*/==-10'd323+xpc10nz) || (4'd12/*MS*/==-10'd322+xpc10nz) || (4'd12/*MS*/==-10'd321+xpc10nz) || (4'd12/*MS*/==
              -10'd320+xpc10nz) || (4'd12/*MS*/==-10'd319+xpc10nz) || (4'd12/*MS*/==-10'd318+xpc10nz) || (4'd12/*MS*/==-10'd314+xpc10nz
              ) || (4'd12/*MS*/==-10'd289+xpc10nz) || (4'd12/*MS*/==-10'd287+xpc10nz) || (4'd12/*MS*/==-10'd285+xpc10nz) || (4'd12/*MS*/==
              -10'd284+xpc10nz) || (4'd12/*MS*/==-10'd259+xpc10nz) || (4'd12/*MS*/==-10'd258+xpc10nz) || (4'd12/*MS*/==-10'd257+xpc10nz
              ) || (4'd12/*MS*/==-9'd255+xpc10nz) || (4'd12/*MS*/==-9'd254+xpc10nz) || (4'd12/*MS*/==-9'd253+xpc10nz) || (4'd12/*MS*/==
              -9'd252+xpc10nz) || (4'd12/*MS*/==-9'd251+xpc10nz) || (4'd12/*MS*/==-9'd250+xpc10nz) || (4'd12/*MS*/==-9'd249+xpc10nz) || 
              (4'd12/*MS*/==-9'd248+xpc10nz) || (4'd12/*MS*/==-9'd247+xpc10nz) || (4'd12/*MS*/==-9'd246+xpc10nz) || (4'd12/*MS*/==-9'd245
              +xpc10nz) || (4'd12/*MS*/==-9'd244+xpc10nz) || (4'd12/*MS*/==-9'd242+xpc10nz) || (4'd12/*MS*/==-9'd241+xpc10nz) || (4'd12
              /*MS*/==-9'd239+xpc10nz) || (4'd12/*MS*/==-9'd238+xpc10nz) || (4'd12/*MS*/==-9'd236+xpc10nz) || (4'd12/*MS*/==-9'd171+xpc10nz
              ) || (4'd12/*MS*/==-8'd106+xpc10nz) || (4'd12/*MS*/==-8'd105+xpc10nz) || (4'd12/*MS*/==-8'd104+xpc10nz) || (4'd12/*MS*/==
              -8'd103+xpc10nz) || (4'd12/*MS*/==-8'd102+xpc10nz) || (4'd12/*MS*/==-8'd101+xpc10nz) || (4'd12/*MS*/==-8'd100+xpc10nz) || 
              (4'd12/*MS*/==-8'd99+xpc10nz) || (4'd12/*MS*/==-8'd98+xpc10nz) || (4'd12/*MS*/==-8'd97+xpc10nz) || (4'd12/*MS*/==-8'd96
              +xpc10nz) || (4'd12/*MS*/==-8'd95+xpc10nz) || (4'd12/*MS*/==-8'd94+xpc10nz) || (4'd12/*MS*/==-8'd93+xpc10nz) || (4'd12/*MS*/==
              -8'd92+xpc10nz) || (4'd12/*MS*/==-8'd91+xpc10nz) || (4'd12/*MS*/==-8'd90+xpc10nz) || (4'd12/*MS*/==-8'd89+xpc10nz) || (4'd12
              /*MS*/==-8'd88+xpc10nz) || (4'd12/*MS*/==-8'd87+xpc10nz) || (4'd12/*MS*/==-8'd86+xpc10nz) || (4'd12/*MS*/==-8'd85+xpc10nz
              ) || (4'd12/*MS*/==-8'd84+xpc10nz) || (4'd12/*MS*/==-8'd83+xpc10nz) || (4'd12/*MS*/==-8'd82+xpc10nz) || (4'd12/*MS*/==-8'd65
              +xpc10nz) || (4'd12/*MS*/==-8'd64+xpc10nz) || (4'd12/*MS*/==-7'd59+xpc10nz) || (4'd12/*MS*/==-7'd50+xpc10nz) || (4'd12/*MS*/==
              -7'd37+xpc10nz) || (4'd12/*MS*/==-6'd20+xpc10nz) || (4'd12/*MS*/==-6'd19+xpc10nz) || (4'd12/*MS*/==-6'd18+xpc10nz) || (4'd12
              /*MS*/==-6'd17+xpc10nz) || (4'd12/*MS*/==-6'd16+xpc10nz) || (4'd12/*MS*/==-5'd15+xpc10nz) || (4'd12/*MS*/==-5'd14+xpc10nz
              ) || (4'd12/*MS*/==-5'd13+xpc10nz) || (4'd12/*MS*/==-5'd12+xpc10nz) || (4'd12/*MS*/==-5'd11+xpc10nz) || (4'd12/*MS*/==-5'd10
              +xpc10nz) || (4'd12/*MS*/==-5'd9+xpc10nz) || (4'd12/*MS*/==-5'd8+xpc10nz) || (4'd12/*MS*/==-4'd7+xpc10nz) || (4'd12/*MS*/==
              -4'd6+xpc10nz) || (4'd12/*MS*/==-4'd5+xpc10nz) || (4'd12/*MS*/==-4'd4+xpc10nz) || (4'd12/*MS*/==-3'd3+xpc10nz) || (4'd12
              /*MS*/==-3'd2+xpc10nz) || (4'd12/*MS*/==-2'd1+xpc10nz) || (xpc10nz==4'd12/*US*/)) && !xpc10_clear && !xpc10_stall;

               xpc10_trk11 <= ((4'd11/*MS*/==-11'd609+xpc10nz) || (4'd11/*MS*/==-11'd599+xpc10nz) || (4'd11/*MS*/==-11'd588+xpc10nz) || 
              (4'd11/*MS*/==-11'd576+xpc10nz) || (4'd11/*MS*/==-11'd571+xpc10nz) || (4'd11/*MS*/==-11'd565+xpc10nz) || (4'd11/*MS*/==
              -11'd558+xpc10nz) || (4'd11/*MS*/==-11'd550+xpc10nz) || (4'd11/*MS*/==-11'd549+xpc10nz) || (4'd11/*MS*/==-11'd547+xpc10nz
              ) || (4'd11/*MS*/==-11'd544+xpc10nz) || (4'd11/*MS*/==-11'd540+xpc10nz) || (4'd11/*MS*/==-11'd539+xpc10nz) || (4'd11/*MS*/==
              -11'd537+xpc10nz) || (4'd11/*MS*/==-11'd534+xpc10nz) || (4'd11/*MS*/==-11'd532+xpc10nz) || (4'd11/*MS*/==-11'd528+xpc10nz
              ) || (4'd11/*MS*/==-10'd503+xpc10nz) || (4'd11/*MS*/==-10'd502+xpc10nz) || (4'd11/*MS*/==-10'd472+xpc10nz) || (4'd11/*MS*/==
              -10'd407+xpc10nz) || (4'd11/*MS*/==-10'd342+xpc10nz) || (4'd11/*MS*/==-10'd341+xpc10nz) || (4'd11/*MS*/==-10'd340+xpc10nz
              ) || (4'd11/*MS*/==-10'd338+xpc10nz) || (4'd11/*MS*/==-10'd335+xpc10nz) || (4'd11/*MS*/==-10'd334+xpc10nz) || (4'd11/*MS*/==
              -10'd330+xpc10nz) || (4'd11/*MS*/==-10'd329+xpc10nz) || (4'd11/*MS*/==-10'd327+xpc10nz) || (4'd11/*MS*/==-10'd324+xpc10nz
              ) || (4'd11/*MS*/==-10'd323+xpc10nz) || (4'd11/*MS*/==-10'd322+xpc10nz) || (4'd11/*MS*/==-10'd321+xpc10nz) || (4'd11/*MS*/==
              -10'd320+xpc10nz) || (4'd11/*MS*/==-10'd319+xpc10nz) || (4'd11/*MS*/==-10'd318+xpc10nz) || (4'd11/*MS*/==-10'd314+xpc10nz
              ) || (4'd11/*MS*/==-10'd289+xpc10nz) || (4'd11/*MS*/==-10'd287+xpc10nz) || (4'd11/*MS*/==-10'd285+xpc10nz) || (4'd11/*MS*/==
              -10'd284+xpc10nz) || (4'd11/*MS*/==-10'd259+xpc10nz) || (4'd11/*MS*/==-10'd258+xpc10nz) || (4'd11/*MS*/==-10'd257+xpc10nz
              ) || (4'd11/*MS*/==-9'd255+xpc10nz) || (4'd11/*MS*/==-9'd254+xpc10nz) || (4'd11/*MS*/==-9'd253+xpc10nz) || (4'd11/*MS*/==
              -9'd252+xpc10nz) || (4'd11/*MS*/==-9'd251+xpc10nz) || (4'd11/*MS*/==-9'd250+xpc10nz) || (4'd11/*MS*/==-9'd249+xpc10nz) || 
              (4'd11/*MS*/==-9'd248+xpc10nz) || (4'd11/*MS*/==-9'd247+xpc10nz) || (4'd11/*MS*/==-9'd246+xpc10nz) || (4'd11/*MS*/==-9'd245
              +xpc10nz) || (4'd11/*MS*/==-9'd244+xpc10nz) || (4'd11/*MS*/==-9'd242+xpc10nz) || (4'd11/*MS*/==-9'd241+xpc10nz) || (4'd11
              /*MS*/==-9'd239+xpc10nz) || (4'd11/*MS*/==-9'd238+xpc10nz) || (4'd11/*MS*/==-9'd236+xpc10nz) || (4'd11/*MS*/==-9'd171+xpc10nz
              ) || (4'd11/*MS*/==-8'd106+xpc10nz) || (4'd11/*MS*/==-8'd105+xpc10nz) || (4'd11/*MS*/==-8'd104+xpc10nz) || (4'd11/*MS*/==
              -8'd103+xpc10nz) || (4'd11/*MS*/==-8'd102+xpc10nz) || (4'd11/*MS*/==-8'd101+xpc10nz) || (4'd11/*MS*/==-8'd100+xpc10nz) || 
              (4'd11/*MS*/==-8'd99+xpc10nz) || (4'd11/*MS*/==-8'd98+xpc10nz) || (4'd11/*MS*/==-8'd97+xpc10nz) || (4'd11/*MS*/==-8'd96
              +xpc10nz) || (4'd11/*MS*/==-8'd95+xpc10nz) || (4'd11/*MS*/==-8'd94+xpc10nz) || (4'd11/*MS*/==-8'd93+xpc10nz) || (4'd11/*MS*/==
              -8'd92+xpc10nz) || (4'd11/*MS*/==-8'd91+xpc10nz) || (4'd11/*MS*/==-8'd90+xpc10nz) || (4'd11/*MS*/==-8'd89+xpc10nz) || (4'd11
              /*MS*/==-8'd88+xpc10nz) || (4'd11/*MS*/==-8'd87+xpc10nz) || (4'd11/*MS*/==-8'd86+xpc10nz) || (4'd11/*MS*/==-8'd85+xpc10nz
              ) || (4'd11/*MS*/==-8'd84+xpc10nz) || (4'd11/*MS*/==-8'd83+xpc10nz) || (4'd11/*MS*/==-8'd82+xpc10nz) || (4'd11/*MS*/==-8'd65
              +xpc10nz) || (4'd11/*MS*/==-8'd64+xpc10nz) || (4'd11/*MS*/==-7'd59+xpc10nz) || (4'd11/*MS*/==-7'd50+xpc10nz) || (4'd11/*MS*/==
              -7'd37+xpc10nz) || (4'd11/*MS*/==-6'd20+xpc10nz) || (4'd11/*MS*/==-6'd19+xpc10nz) || (4'd11/*MS*/==-6'd18+xpc10nz) || (4'd11
              /*MS*/==-6'd17+xpc10nz) || (4'd11/*MS*/==-6'd16+xpc10nz) || (4'd11/*MS*/==-5'd15+xpc10nz) || (4'd11/*MS*/==-5'd14+xpc10nz
              ) || (4'd11/*MS*/==-5'd13+xpc10nz) || (4'd11/*MS*/==-5'd12+xpc10nz) || (4'd11/*MS*/==-5'd11+xpc10nz) || (4'd11/*MS*/==-5'd10
              +xpc10nz) || (4'd11/*MS*/==-5'd9+xpc10nz) || (4'd11/*MS*/==-5'd8+xpc10nz) || (4'd11/*MS*/==-4'd7+xpc10nz) || (4'd11/*MS*/==
              -4'd6+xpc10nz) || (4'd11/*MS*/==-4'd5+xpc10nz) || (4'd11/*MS*/==-4'd4+xpc10nz) || (4'd11/*MS*/==-3'd3+xpc10nz) || (4'd11
              /*MS*/==-3'd2+xpc10nz) || (4'd11/*MS*/==-2'd1+xpc10nz) || (xpc10nz==4'd11/*US*/)) && !xpc10_clear && !xpc10_stall;

               xpc10_trk10 <= ((4'd10/*MS*/==-11'd609+xpc10nz) || (4'd10/*MS*/==-11'd599+xpc10nz) || (4'd10/*MS*/==-11'd588+xpc10nz) || 
              (4'd10/*MS*/==-11'd576+xpc10nz) || (4'd10/*MS*/==-11'd571+xpc10nz) || (4'd10/*MS*/==-11'd565+xpc10nz) || (4'd10/*MS*/==
              -11'd558+xpc10nz) || (4'd10/*MS*/==-11'd550+xpc10nz) || (4'd10/*MS*/==-11'd549+xpc10nz) || (4'd10/*MS*/==-11'd547+xpc10nz
              ) || (4'd10/*MS*/==-11'd544+xpc10nz) || (4'd10/*MS*/==-11'd540+xpc10nz) || (4'd10/*MS*/==-11'd539+xpc10nz) || (4'd10/*MS*/==
              -11'd537+xpc10nz) || (4'd10/*MS*/==-11'd534+xpc10nz) || (4'd10/*MS*/==-11'd532+xpc10nz) || (4'd10/*MS*/==-11'd528+xpc10nz
              ) || (4'd10/*MS*/==-10'd503+xpc10nz) || (4'd10/*MS*/==-10'd502+xpc10nz) || (4'd10/*MS*/==-10'd472+xpc10nz) || (4'd10/*MS*/==
              -10'd407+xpc10nz) || (4'd10/*MS*/==-10'd342+xpc10nz) || (4'd10/*MS*/==-10'd341+xpc10nz) || (4'd10/*MS*/==-10'd340+xpc10nz
              ) || (4'd10/*MS*/==-10'd338+xpc10nz) || (4'd10/*MS*/==-10'd335+xpc10nz) || (4'd10/*MS*/==-10'd334+xpc10nz) || (4'd10/*MS*/==
              -10'd330+xpc10nz) || (4'd10/*MS*/==-10'd329+xpc10nz) || (4'd10/*MS*/==-10'd327+xpc10nz) || (4'd10/*MS*/==-10'd324+xpc10nz
              ) || (4'd10/*MS*/==-10'd323+xpc10nz) || (4'd10/*MS*/==-10'd322+xpc10nz) || (4'd10/*MS*/==-10'd321+xpc10nz) || (4'd10/*MS*/==
              -10'd320+xpc10nz) || (4'd10/*MS*/==-10'd319+xpc10nz) || (4'd10/*MS*/==-10'd318+xpc10nz) || (4'd10/*MS*/==-10'd314+xpc10nz
              ) || (4'd10/*MS*/==-10'd289+xpc10nz) || (4'd10/*MS*/==-10'd287+xpc10nz) || (4'd10/*MS*/==-10'd285+xpc10nz) || (4'd10/*MS*/==
              -10'd284+xpc10nz) || (4'd10/*MS*/==-10'd259+xpc10nz) || (4'd10/*MS*/==-10'd258+xpc10nz) || (4'd10/*MS*/==-10'd257+xpc10nz
              ) || (4'd10/*MS*/==-9'd255+xpc10nz) || (4'd10/*MS*/==-9'd254+xpc10nz) || (4'd10/*MS*/==-9'd253+xpc10nz) || (4'd10/*MS*/==
              -9'd252+xpc10nz) || (4'd10/*MS*/==-9'd251+xpc10nz) || (4'd10/*MS*/==-9'd250+xpc10nz) || (4'd10/*MS*/==-9'd249+xpc10nz) || 
              (4'd10/*MS*/==-9'd248+xpc10nz) || (4'd10/*MS*/==-9'd247+xpc10nz) || (4'd10/*MS*/==-9'd246+xpc10nz) || (4'd10/*MS*/==-9'd245
              +xpc10nz) || (4'd10/*MS*/==-9'd244+xpc10nz) || (4'd10/*MS*/==-9'd242+xpc10nz) || (4'd10/*MS*/==-9'd241+xpc10nz) || (4'd10
              /*MS*/==-9'd239+xpc10nz) || (4'd10/*MS*/==-9'd238+xpc10nz) || (4'd10/*MS*/==-9'd236+xpc10nz) || (4'd10/*MS*/==-9'd171+xpc10nz
              ) || (4'd10/*MS*/==-8'd106+xpc10nz) || (4'd10/*MS*/==-8'd105+xpc10nz) || (4'd10/*MS*/==-8'd104+xpc10nz) || (4'd10/*MS*/==
              -8'd103+xpc10nz) || (4'd10/*MS*/==-8'd102+xpc10nz) || (4'd10/*MS*/==-8'd101+xpc10nz) || (4'd10/*MS*/==-8'd100+xpc10nz) || 
              (4'd10/*MS*/==-8'd99+xpc10nz) || (4'd10/*MS*/==-8'd98+xpc10nz) || (4'd10/*MS*/==-8'd97+xpc10nz) || (4'd10/*MS*/==-8'd96
              +xpc10nz) || (4'd10/*MS*/==-8'd95+xpc10nz) || (4'd10/*MS*/==-8'd94+xpc10nz) || (4'd10/*MS*/==-8'd93+xpc10nz) || (4'd10/*MS*/==
              -8'd92+xpc10nz) || (4'd10/*MS*/==-8'd91+xpc10nz) || (4'd10/*MS*/==-8'd90+xpc10nz) || (4'd10/*MS*/==-8'd89+xpc10nz) || (4'd10
              /*MS*/==-8'd88+xpc10nz) || (4'd10/*MS*/==-8'd87+xpc10nz) || (4'd10/*MS*/==-8'd86+xpc10nz) || (4'd10/*MS*/==-8'd85+xpc10nz
              ) || (4'd10/*MS*/==-8'd84+xpc10nz) || (4'd10/*MS*/==-8'd83+xpc10nz) || (4'd10/*MS*/==-8'd82+xpc10nz) || (4'd10/*MS*/==-8'd65
              +xpc10nz) || (4'd10/*MS*/==-8'd64+xpc10nz) || (4'd10/*MS*/==-7'd59+xpc10nz) || (4'd10/*MS*/==-7'd50+xpc10nz) || (4'd10/*MS*/==
              -7'd37+xpc10nz) || (4'd10/*MS*/==-6'd20+xpc10nz) || (4'd10/*MS*/==-6'd19+xpc10nz) || (4'd10/*MS*/==-6'd18+xpc10nz) || (4'd10
              /*MS*/==-6'd17+xpc10nz) || (4'd10/*MS*/==-6'd16+xpc10nz) || (4'd10/*MS*/==-5'd15+xpc10nz) || (4'd10/*MS*/==-5'd14+xpc10nz
              ) || (4'd10/*MS*/==-5'd13+xpc10nz) || (4'd10/*MS*/==-5'd12+xpc10nz) || (4'd10/*MS*/==-5'd11+xpc10nz) || (4'd10/*MS*/==-5'd10
              +xpc10nz) || (4'd10/*MS*/==-5'd9+xpc10nz) || (4'd10/*MS*/==-5'd8+xpc10nz) || (4'd10/*MS*/==-4'd7+xpc10nz) || (4'd10/*MS*/==
              -4'd6+xpc10nz) || (4'd10/*MS*/==-4'd5+xpc10nz) || (4'd10/*MS*/==-4'd4+xpc10nz) || (4'd10/*MS*/==-3'd3+xpc10nz) || (4'd10
              /*MS*/==-3'd2+xpc10nz) || (4'd10/*MS*/==-2'd1+xpc10nz) || (xpc10nz==4'd10/*US*/)) && !xpc10_clear && !xpc10_stall;

               xpc10_trk9 <= ((4'd9/*MS*/==-11'd609+xpc10nz) || (4'd9/*MS*/==-11'd599+xpc10nz) || (4'd9/*MS*/==-11'd588+xpc10nz) || (4'd9
              /*MS*/==-11'd576+xpc10nz) || (4'd9/*MS*/==-11'd571+xpc10nz) || (4'd9/*MS*/==-11'd565+xpc10nz) || (4'd9/*MS*/==-11'd558+
              xpc10nz) || (4'd9/*MS*/==-11'd550+xpc10nz) || (4'd9/*MS*/==-11'd549+xpc10nz) || (4'd9/*MS*/==-11'd547+xpc10nz) || (4'd9
              /*MS*/==-11'd544+xpc10nz) || (4'd9/*MS*/==-11'd540+xpc10nz) || (4'd9/*MS*/==-11'd539+xpc10nz) || (4'd9/*MS*/==-11'd537+
              xpc10nz) || (4'd9/*MS*/==-11'd534+xpc10nz) || (4'd9/*MS*/==-11'd532+xpc10nz) || (4'd9/*MS*/==-11'd528+xpc10nz) || (4'd9
              /*MS*/==-10'd503+xpc10nz) || (4'd9/*MS*/==-10'd502+xpc10nz) || (4'd9/*MS*/==-10'd472+xpc10nz) || (4'd9/*MS*/==-10'd407+
              xpc10nz) || (4'd9/*MS*/==-10'd342+xpc10nz) || (4'd9/*MS*/==-10'd341+xpc10nz) || (4'd9/*MS*/==-10'd340+xpc10nz) || (4'd9
              /*MS*/==-10'd338+xpc10nz) || (4'd9/*MS*/==-10'd335+xpc10nz) || (4'd9/*MS*/==-10'd334+xpc10nz) || (4'd9/*MS*/==-10'd330+
              xpc10nz) || (4'd9/*MS*/==-10'd329+xpc10nz) || (4'd9/*MS*/==-10'd327+xpc10nz) || (4'd9/*MS*/==-10'd324+xpc10nz) || (4'd9
              /*MS*/==-10'd323+xpc10nz) || (4'd9/*MS*/==-10'd322+xpc10nz) || (4'd9/*MS*/==-10'd321+xpc10nz) || (4'd9/*MS*/==-10'd320+
              xpc10nz) || (4'd9/*MS*/==-10'd319+xpc10nz) || (4'd9/*MS*/==-10'd318+xpc10nz) || (4'd9/*MS*/==-10'd314+xpc10nz) || (4'd9
              /*MS*/==-10'd289+xpc10nz) || (4'd9/*MS*/==-10'd287+xpc10nz) || (4'd9/*MS*/==-10'd285+xpc10nz) || (4'd9/*MS*/==-10'd284+
              xpc10nz) || (4'd9/*MS*/==-10'd259+xpc10nz) || (4'd9/*MS*/==-10'd258+xpc10nz) || (4'd9/*MS*/==-10'd257+xpc10nz) || (4'd9
              /*MS*/==-9'd255+xpc10nz) || (4'd9/*MS*/==-9'd254+xpc10nz) || (4'd9/*MS*/==-9'd253+xpc10nz) || (4'd9/*MS*/==-9'd252+xpc10nz
              ) || (4'd9/*MS*/==-9'd251+xpc10nz) || (4'd9/*MS*/==-9'd250+xpc10nz) || (4'd9/*MS*/==-9'd249+xpc10nz) || (4'd9/*MS*/==-9'd248
              +xpc10nz) || (4'd9/*MS*/==-9'd247+xpc10nz) || (4'd9/*MS*/==-9'd246+xpc10nz) || (4'd9/*MS*/==-9'd245+xpc10nz) || (4'd9/*MS*/==
              -9'd244+xpc10nz) || (4'd9/*MS*/==-9'd242+xpc10nz) || (4'd9/*MS*/==-9'd241+xpc10nz) || (4'd9/*MS*/==-9'd239+xpc10nz) || 
              (4'd9/*MS*/==-9'd238+xpc10nz) || (4'd9/*MS*/==-9'd236+xpc10nz) || (4'd9/*MS*/==-9'd171+xpc10nz) || (4'd9/*MS*/==-8'd106
              +xpc10nz) || (4'd9/*MS*/==-8'd105+xpc10nz) || (4'd9/*MS*/==-8'd104+xpc10nz) || (4'd9/*MS*/==-8'd103+xpc10nz) || (4'd9/*MS*/==
              -8'd102+xpc10nz) || (4'd9/*MS*/==-8'd101+xpc10nz) || (4'd9/*MS*/==-8'd100+xpc10nz) || (4'd9/*MS*/==-8'd99+xpc10nz) || (4'd9
              /*MS*/==-8'd98+xpc10nz) || (4'd9/*MS*/==-8'd97+xpc10nz) || (4'd9/*MS*/==-8'd96+xpc10nz) || (4'd9/*MS*/==-8'd95+xpc10nz) || 
              (4'd9/*MS*/==-8'd94+xpc10nz) || (4'd9/*MS*/==-8'd93+xpc10nz) || (4'd9/*MS*/==-8'd92+xpc10nz) || (4'd9/*MS*/==-8'd91+xpc10nz
              ) || (4'd9/*MS*/==-8'd90+xpc10nz) || (4'd9/*MS*/==-8'd89+xpc10nz) || (4'd9/*MS*/==-8'd88+xpc10nz) || (4'd9/*MS*/==-8'd87
              +xpc10nz) || (4'd9/*MS*/==-8'd86+xpc10nz) || (4'd9/*MS*/==-8'd85+xpc10nz) || (4'd9/*MS*/==-8'd84+xpc10nz) || (4'd9/*MS*/==
              -8'd83+xpc10nz) || (4'd9/*MS*/==-8'd82+xpc10nz) || (4'd9/*MS*/==-8'd65+xpc10nz) || (4'd9/*MS*/==-8'd64+xpc10nz) || (4'd9
              /*MS*/==-7'd59+xpc10nz) || (4'd9/*MS*/==-7'd50+xpc10nz) || (4'd9/*MS*/==-7'd37+xpc10nz) || (4'd9/*MS*/==-6'd20+xpc10nz) || 
              (4'd9/*MS*/==-6'd19+xpc10nz) || (4'd9/*MS*/==-6'd18+xpc10nz) || (4'd9/*MS*/==-6'd17+xpc10nz) || (4'd9/*MS*/==-6'd16+xpc10nz
              ) || (4'd9/*MS*/==-5'd15+xpc10nz) || (4'd9/*MS*/==-5'd14+xpc10nz) || (4'd9/*MS*/==-5'd13+xpc10nz) || (4'd9/*MS*/==-5'd12
              +xpc10nz) || (4'd9/*MS*/==-5'd11+xpc10nz) || (4'd9/*MS*/==-5'd10+xpc10nz) || (4'd9/*MS*/==-5'd9+xpc10nz) || (4'd9/*MS*/==
              -5'd8+xpc10nz) || (4'd9/*MS*/==-4'd7+xpc10nz) || (4'd9/*MS*/==-4'd6+xpc10nz) || (4'd9/*MS*/==-4'd5+xpc10nz) || (4'd9/*MS*/==
              -4'd4+xpc10nz) || (4'd9/*MS*/==-3'd3+xpc10nz) || (4'd9/*MS*/==-3'd2+xpc10nz) || (4'd9/*MS*/==-2'd1+xpc10nz) || (xpc10nz
              ==4'd9/*US*/)) && !xpc10_clear && !xpc10_stall;

               xpc10_trk8 <= ((4'd8/*MS*/==-11'd609+xpc10nz) || (4'd8/*MS*/==-11'd599+xpc10nz) || (4'd8/*MS*/==-11'd588+xpc10nz) || (4'd8
              /*MS*/==-11'd576+xpc10nz) || (4'd8/*MS*/==-11'd571+xpc10nz) || (4'd8/*MS*/==-11'd565+xpc10nz) || (4'd8/*MS*/==-11'd558+
              xpc10nz) || (4'd8/*MS*/==-11'd550+xpc10nz) || (4'd8/*MS*/==-11'd549+xpc10nz) || (4'd8/*MS*/==-11'd547+xpc10nz) || (4'd8
              /*MS*/==-11'd544+xpc10nz) || (4'd8/*MS*/==-11'd540+xpc10nz) || (4'd8/*MS*/==-11'd539+xpc10nz) || (4'd8/*MS*/==-11'd537+
              xpc10nz) || (4'd8/*MS*/==-11'd534+xpc10nz) || (4'd8/*MS*/==-11'd532+xpc10nz) || (4'd8/*MS*/==-11'd528+xpc10nz) || (4'd8
              /*MS*/==-10'd503+xpc10nz) || (4'd8/*MS*/==-10'd502+xpc10nz) || (4'd8/*MS*/==-10'd472+xpc10nz) || (4'd8/*MS*/==-10'd407+
              xpc10nz) || (4'd8/*MS*/==-10'd342+xpc10nz) || (4'd8/*MS*/==-10'd341+xpc10nz) || (4'd8/*MS*/==-10'd340+xpc10nz) || (4'd8
              /*MS*/==-10'd338+xpc10nz) || (4'd8/*MS*/==-10'd335+xpc10nz) || (4'd8/*MS*/==-10'd334+xpc10nz) || (4'd8/*MS*/==-10'd330+
              xpc10nz) || (4'd8/*MS*/==-10'd329+xpc10nz) || (4'd8/*MS*/==-10'd327+xpc10nz) || (4'd8/*MS*/==-10'd324+xpc10nz) || (4'd8
              /*MS*/==-10'd323+xpc10nz) || (4'd8/*MS*/==-10'd322+xpc10nz) || (4'd8/*MS*/==-10'd321+xpc10nz) || (4'd8/*MS*/==-10'd320+
              xpc10nz) || (4'd8/*MS*/==-10'd319+xpc10nz) || (4'd8/*MS*/==-10'd318+xpc10nz) || (4'd8/*MS*/==-10'd314+xpc10nz) || (4'd8
              /*MS*/==-10'd289+xpc10nz) || (4'd8/*MS*/==-10'd287+xpc10nz) || (4'd8/*MS*/==-10'd285+xpc10nz) || (4'd8/*MS*/==-10'd284+
              xpc10nz) || (4'd8/*MS*/==-10'd259+xpc10nz) || (4'd8/*MS*/==-10'd258+xpc10nz) || (4'd8/*MS*/==-10'd257+xpc10nz) || (4'd8
              /*MS*/==-9'd255+xpc10nz) || (4'd8/*MS*/==-9'd254+xpc10nz) || (4'd8/*MS*/==-9'd253+xpc10nz) || (4'd8/*MS*/==-9'd252+xpc10nz
              ) || (4'd8/*MS*/==-9'd251+xpc10nz) || (4'd8/*MS*/==-9'd250+xpc10nz) || (4'd8/*MS*/==-9'd249+xpc10nz) || (4'd8/*MS*/==-9'd248
              +xpc10nz) || (4'd8/*MS*/==-9'd247+xpc10nz) || (4'd8/*MS*/==-9'd246+xpc10nz) || (4'd8/*MS*/==-9'd245+xpc10nz) || (4'd8/*MS*/==
              -9'd244+xpc10nz) || (4'd8/*MS*/==-9'd242+xpc10nz) || (4'd8/*MS*/==-9'd241+xpc10nz) || (4'd8/*MS*/==-9'd239+xpc10nz) || 
              (4'd8/*MS*/==-9'd238+xpc10nz) || (4'd8/*MS*/==-9'd236+xpc10nz) || (4'd8/*MS*/==-9'd171+xpc10nz) || (4'd8/*MS*/==-8'd106
              +xpc10nz) || (4'd8/*MS*/==-8'd105+xpc10nz) || (4'd8/*MS*/==-8'd104+xpc10nz) || (4'd8/*MS*/==-8'd103+xpc10nz) || (4'd8/*MS*/==
              -8'd102+xpc10nz) || (4'd8/*MS*/==-8'd101+xpc10nz) || (4'd8/*MS*/==-8'd100+xpc10nz) || (4'd8/*MS*/==-8'd99+xpc10nz) || (4'd8
              /*MS*/==-8'd98+xpc10nz) || (4'd8/*MS*/==-8'd97+xpc10nz) || (4'd8/*MS*/==-8'd96+xpc10nz) || (4'd8/*MS*/==-8'd95+xpc10nz) || 
              (4'd8/*MS*/==-8'd94+xpc10nz) || (4'd8/*MS*/==-8'd93+xpc10nz) || (4'd8/*MS*/==-8'd92+xpc10nz) || (4'd8/*MS*/==-8'd91+xpc10nz
              ) || (4'd8/*MS*/==-8'd90+xpc10nz) || (4'd8/*MS*/==-8'd89+xpc10nz) || (4'd8/*MS*/==-8'd88+xpc10nz) || (4'd8/*MS*/==-8'd87
              +xpc10nz) || (4'd8/*MS*/==-8'd86+xpc10nz) || (4'd8/*MS*/==-8'd85+xpc10nz) || (4'd8/*MS*/==-8'd84+xpc10nz) || (4'd8/*MS*/==
              -8'd83+xpc10nz) || (4'd8/*MS*/==-8'd82+xpc10nz) || (4'd8/*MS*/==-8'd65+xpc10nz) || (4'd8/*MS*/==-8'd64+xpc10nz) || (4'd8
              /*MS*/==-7'd59+xpc10nz) || (4'd8/*MS*/==-7'd50+xpc10nz) || (4'd8/*MS*/==-7'd37+xpc10nz) || (4'd8/*MS*/==-6'd20+xpc10nz) || 
              (4'd8/*MS*/==-6'd19+xpc10nz) || (4'd8/*MS*/==-6'd18+xpc10nz) || (4'd8/*MS*/==-6'd17+xpc10nz) || (4'd8/*MS*/==-6'd16+xpc10nz
              ) || (4'd8/*MS*/==-5'd15+xpc10nz) || (4'd8/*MS*/==-5'd14+xpc10nz) || (4'd8/*MS*/==-5'd13+xpc10nz) || (4'd8/*MS*/==-5'd12
              +xpc10nz) || (4'd8/*MS*/==-5'd11+xpc10nz) || (4'd8/*MS*/==-5'd10+xpc10nz) || (4'd8/*MS*/==-5'd9+xpc10nz) || (4'd8/*MS*/==
              -5'd8+xpc10nz) || (4'd8/*MS*/==-4'd7+xpc10nz) || (4'd8/*MS*/==-4'd6+xpc10nz) || (4'd8/*MS*/==-4'd5+xpc10nz) || (4'd8/*MS*/==
              -4'd4+xpc10nz) || (4'd8/*MS*/==-3'd3+xpc10nz) || (4'd8/*MS*/==-3'd2+xpc10nz) || (4'd8/*MS*/==-2'd1+xpc10nz) || (xpc10nz
              ==4'd8/*US*/)) && !xpc10_clear && !xpc10_stall;

               xpc10_trk7 <= ((3'd7/*MS*/==-11'd609+xpc10nz) || (3'd7/*MS*/==-11'd599+xpc10nz) || (3'd7/*MS*/==-11'd588+xpc10nz) || (3'd7
              /*MS*/==-11'd576+xpc10nz) || (3'd7/*MS*/==-11'd571+xpc10nz) || (3'd7/*MS*/==-11'd565+xpc10nz) || (3'd7/*MS*/==-11'd558+
              xpc10nz) || (3'd7/*MS*/==-11'd550+xpc10nz) || (3'd7/*MS*/==-11'd549+xpc10nz) || (3'd7/*MS*/==-11'd547+xpc10nz) || (3'd7
              /*MS*/==-11'd544+xpc10nz) || (3'd7/*MS*/==-11'd540+xpc10nz) || (3'd7/*MS*/==-11'd539+xpc10nz) || (3'd7/*MS*/==-11'd537+
              xpc10nz) || (3'd7/*MS*/==-11'd534+xpc10nz) || (3'd7/*MS*/==-11'd532+xpc10nz) || (3'd7/*MS*/==-11'd528+xpc10nz) || (3'd7
              /*MS*/==-10'd503+xpc10nz) || (3'd7/*MS*/==-10'd502+xpc10nz) || (3'd7/*MS*/==-10'd472+xpc10nz) || (3'd7/*MS*/==-10'd407+
              xpc10nz) || (3'd7/*MS*/==-10'd342+xpc10nz) || (3'd7/*MS*/==-10'd341+xpc10nz) || (3'd7/*MS*/==-10'd340+xpc10nz) || (3'd7
              /*MS*/==-10'd338+xpc10nz) || (3'd7/*MS*/==-10'd335+xpc10nz) || (3'd7/*MS*/==-10'd334+xpc10nz) || (3'd7/*MS*/==-10'd330+
              xpc10nz) || (3'd7/*MS*/==-10'd329+xpc10nz) || (3'd7/*MS*/==-10'd327+xpc10nz) || (3'd7/*MS*/==-10'd324+xpc10nz) || (3'd7
              /*MS*/==-10'd323+xpc10nz) || (3'd7/*MS*/==-10'd322+xpc10nz) || (3'd7/*MS*/==-10'd321+xpc10nz) || (3'd7/*MS*/==-10'd320+
              xpc10nz) || (3'd7/*MS*/==-10'd319+xpc10nz) || (3'd7/*MS*/==-10'd318+xpc10nz) || (3'd7/*MS*/==-10'd314+xpc10nz) || (3'd7
              /*MS*/==-10'd289+xpc10nz) || (3'd7/*MS*/==-10'd287+xpc10nz) || (3'd7/*MS*/==-10'd285+xpc10nz) || (3'd7/*MS*/==-10'd284+
              xpc10nz) || (3'd7/*MS*/==-10'd259+xpc10nz) || (3'd7/*MS*/==-10'd258+xpc10nz) || (3'd7/*MS*/==-10'd257+xpc10nz) || (3'd7
              /*MS*/==-9'd255+xpc10nz) || (3'd7/*MS*/==-9'd254+xpc10nz) || (3'd7/*MS*/==-9'd253+xpc10nz) || (3'd7/*MS*/==-9'd252+xpc10nz
              ) || (3'd7/*MS*/==-9'd251+xpc10nz) || (3'd7/*MS*/==-9'd250+xpc10nz) || (3'd7/*MS*/==-9'd249+xpc10nz) || (3'd7/*MS*/==-9'd248
              +xpc10nz) || (3'd7/*MS*/==-9'd247+xpc10nz) || (3'd7/*MS*/==-9'd246+xpc10nz) || (3'd7/*MS*/==-9'd245+xpc10nz) || (3'd7/*MS*/==
              -9'd244+xpc10nz) || (3'd7/*MS*/==-9'd242+xpc10nz) || (3'd7/*MS*/==-9'd241+xpc10nz) || (3'd7/*MS*/==-9'd239+xpc10nz) || 
              (3'd7/*MS*/==-9'd238+xpc10nz) || (3'd7/*MS*/==-9'd236+xpc10nz) || (3'd7/*MS*/==-9'd171+xpc10nz) || (3'd7/*MS*/==-8'd106
              +xpc10nz) || (3'd7/*MS*/==-8'd105+xpc10nz) || (3'd7/*MS*/==-8'd104+xpc10nz) || (3'd7/*MS*/==-8'd103+xpc10nz) || (3'd7/*MS*/==
              -8'd102+xpc10nz) || (3'd7/*MS*/==-8'd101+xpc10nz) || (3'd7/*MS*/==-8'd100+xpc10nz) || (3'd7/*MS*/==-8'd99+xpc10nz) || (3'd7
              /*MS*/==-8'd98+xpc10nz) || (3'd7/*MS*/==-8'd97+xpc10nz) || (3'd7/*MS*/==-8'd96+xpc10nz) || (3'd7/*MS*/==-8'd95+xpc10nz) || 
              (3'd7/*MS*/==-8'd94+xpc10nz) || (3'd7/*MS*/==-8'd93+xpc10nz) || (3'd7/*MS*/==-8'd92+xpc10nz) || (3'd7/*MS*/==-8'd91+xpc10nz
              ) || (3'd7/*MS*/==-8'd90+xpc10nz) || (3'd7/*MS*/==-8'd89+xpc10nz) || (3'd7/*MS*/==-8'd88+xpc10nz) || (3'd7/*MS*/==-8'd87
              +xpc10nz) || (3'd7/*MS*/==-8'd86+xpc10nz) || (3'd7/*MS*/==-8'd85+xpc10nz) || (3'd7/*MS*/==-8'd84+xpc10nz) || (3'd7/*MS*/==
              -8'd83+xpc10nz) || (3'd7/*MS*/==-8'd82+xpc10nz) || (3'd7/*MS*/==-8'd65+xpc10nz) || (3'd7/*MS*/==-8'd64+xpc10nz) || (3'd7
              /*MS*/==-7'd59+xpc10nz) || (3'd7/*MS*/==-7'd50+xpc10nz) || (3'd7/*MS*/==-7'd37+xpc10nz) || (3'd7/*MS*/==-6'd20+xpc10nz) || 
              (3'd7/*MS*/==-6'd19+xpc10nz) || (3'd7/*MS*/==-6'd18+xpc10nz) || (3'd7/*MS*/==-6'd17+xpc10nz) || (3'd7/*MS*/==-6'd16+xpc10nz
              ) || (3'd7/*MS*/==-5'd15+xpc10nz) || (3'd7/*MS*/==-5'd14+xpc10nz) || (3'd7/*MS*/==-5'd13+xpc10nz) || (3'd7/*MS*/==-5'd12
              +xpc10nz) || (3'd7/*MS*/==-5'd11+xpc10nz) || (3'd7/*MS*/==-5'd10+xpc10nz) || (3'd7/*MS*/==-5'd9+xpc10nz) || (3'd7/*MS*/==
              -5'd8+xpc10nz) || (3'd7/*MS*/==-4'd7+xpc10nz) || (3'd7/*MS*/==-4'd6+xpc10nz) || (3'd7/*MS*/==-4'd5+xpc10nz) || (3'd7/*MS*/==
              -4'd4+xpc10nz) || (3'd7/*MS*/==-3'd3+xpc10nz) || (3'd7/*MS*/==-3'd2+xpc10nz) || (3'd7/*MS*/==-2'd1+xpc10nz) || (xpc10nz
              ==3'd7/*US*/)) && !xpc10_clear && !xpc10_stall;

               xpc10_trk6 <= ((3'd6/*MS*/==-11'd609+xpc10nz) || (3'd6/*MS*/==-11'd599+xpc10nz) || (3'd6/*MS*/==-11'd588+xpc10nz) || (3'd6
              /*MS*/==-11'd576+xpc10nz) || (3'd6/*MS*/==-11'd571+xpc10nz) || (3'd6/*MS*/==-11'd565+xpc10nz) || (3'd6/*MS*/==-11'd558+
              xpc10nz) || (3'd6/*MS*/==-11'd550+xpc10nz) || (3'd6/*MS*/==-11'd549+xpc10nz) || (3'd6/*MS*/==-11'd547+xpc10nz) || (3'd6
              /*MS*/==-11'd544+xpc10nz) || (3'd6/*MS*/==-11'd540+xpc10nz) || (3'd6/*MS*/==-11'd539+xpc10nz) || (3'd6/*MS*/==-11'd537+
              xpc10nz) || (3'd6/*MS*/==-11'd534+xpc10nz) || (3'd6/*MS*/==-11'd532+xpc10nz) || (3'd6/*MS*/==-11'd528+xpc10nz) || (3'd6
              /*MS*/==-10'd503+xpc10nz) || (3'd6/*MS*/==-10'd502+xpc10nz) || (3'd6/*MS*/==-10'd472+xpc10nz) || (3'd6/*MS*/==-10'd407+
              xpc10nz) || (3'd6/*MS*/==-10'd342+xpc10nz) || (3'd6/*MS*/==-10'd341+xpc10nz) || (3'd6/*MS*/==-10'd340+xpc10nz) || (3'd6
              /*MS*/==-10'd338+xpc10nz) || (3'd6/*MS*/==-10'd335+xpc10nz) || (3'd6/*MS*/==-10'd334+xpc10nz) || (3'd6/*MS*/==-10'd330+
              xpc10nz) || (3'd6/*MS*/==-10'd329+xpc10nz) || (3'd6/*MS*/==-10'd327+xpc10nz) || (3'd6/*MS*/==-10'd324+xpc10nz) || (3'd6
              /*MS*/==-10'd323+xpc10nz) || (3'd6/*MS*/==-10'd322+xpc10nz) || (3'd6/*MS*/==-10'd321+xpc10nz) || (3'd6/*MS*/==-10'd320+
              xpc10nz) || (3'd6/*MS*/==-10'd319+xpc10nz) || (3'd6/*MS*/==-10'd318+xpc10nz) || (3'd6/*MS*/==-10'd314+xpc10nz) || (3'd6
              /*MS*/==-10'd289+xpc10nz) || (3'd6/*MS*/==-10'd287+xpc10nz) || (3'd6/*MS*/==-10'd285+xpc10nz) || (3'd6/*MS*/==-10'd284+
              xpc10nz) || (3'd6/*MS*/==-10'd259+xpc10nz) || (3'd6/*MS*/==-10'd258+xpc10nz) || (3'd6/*MS*/==-10'd257+xpc10nz) || (3'd6
              /*MS*/==-9'd255+xpc10nz) || (3'd6/*MS*/==-9'd254+xpc10nz) || (3'd6/*MS*/==-9'd253+xpc10nz) || (3'd6/*MS*/==-9'd252+xpc10nz
              ) || (3'd6/*MS*/==-9'd251+xpc10nz) || (3'd6/*MS*/==-9'd250+xpc10nz) || (3'd6/*MS*/==-9'd249+xpc10nz) || (3'd6/*MS*/==-9'd248
              +xpc10nz) || (3'd6/*MS*/==-9'd247+xpc10nz) || (3'd6/*MS*/==-9'd246+xpc10nz) || (3'd6/*MS*/==-9'd245+xpc10nz) || (3'd6/*MS*/==
              -9'd244+xpc10nz) || (3'd6/*MS*/==-9'd242+xpc10nz) || (3'd6/*MS*/==-9'd241+xpc10nz) || (3'd6/*MS*/==-9'd239+xpc10nz) || 
              (3'd6/*MS*/==-9'd238+xpc10nz) || (3'd6/*MS*/==-9'd236+xpc10nz) || (3'd6/*MS*/==-9'd171+xpc10nz) || (3'd6/*MS*/==-8'd106
              +xpc10nz) || (3'd6/*MS*/==-8'd105+xpc10nz) || (3'd6/*MS*/==-8'd104+xpc10nz) || (3'd6/*MS*/==-8'd103+xpc10nz) || (3'd6/*MS*/==
              -8'd102+xpc10nz) || (3'd6/*MS*/==-8'd101+xpc10nz) || (3'd6/*MS*/==-8'd100+xpc10nz) || (3'd6/*MS*/==-8'd99+xpc10nz) || (3'd6
              /*MS*/==-8'd98+xpc10nz) || (3'd6/*MS*/==-8'd97+xpc10nz) || (3'd6/*MS*/==-8'd96+xpc10nz) || (3'd6/*MS*/==-8'd95+xpc10nz) || 
              (3'd6/*MS*/==-8'd94+xpc10nz) || (3'd6/*MS*/==-8'd93+xpc10nz) || (3'd6/*MS*/==-8'd92+xpc10nz) || (3'd6/*MS*/==-8'd91+xpc10nz
              ) || (3'd6/*MS*/==-8'd90+xpc10nz) || (3'd6/*MS*/==-8'd89+xpc10nz) || (3'd6/*MS*/==-8'd88+xpc10nz) || (3'd6/*MS*/==-8'd87
              +xpc10nz) || (3'd6/*MS*/==-8'd86+xpc10nz) || (3'd6/*MS*/==-8'd85+xpc10nz) || (3'd6/*MS*/==-8'd84+xpc10nz) || (3'd6/*MS*/==
              -8'd83+xpc10nz) || (3'd6/*MS*/==-8'd82+xpc10nz) || (3'd6/*MS*/==-8'd65+xpc10nz) || (3'd6/*MS*/==-8'd64+xpc10nz) || (3'd6
              /*MS*/==-7'd59+xpc10nz) || (3'd6/*MS*/==-7'd50+xpc10nz) || (3'd6/*MS*/==-7'd37+xpc10nz) || (3'd6/*MS*/==-6'd20+xpc10nz) || 
              (3'd6/*MS*/==-6'd19+xpc10nz) || (3'd6/*MS*/==-6'd18+xpc10nz) || (3'd6/*MS*/==-6'd17+xpc10nz) || (3'd6/*MS*/==-6'd16+xpc10nz
              ) || (3'd6/*MS*/==-5'd15+xpc10nz) || (3'd6/*MS*/==-5'd14+xpc10nz) || (3'd6/*MS*/==-5'd13+xpc10nz) || (3'd6/*MS*/==-5'd12
              +xpc10nz) || (3'd6/*MS*/==-5'd11+xpc10nz) || (3'd6/*MS*/==-5'd10+xpc10nz) || (3'd6/*MS*/==-5'd9+xpc10nz) || (3'd6/*MS*/==
              -5'd8+xpc10nz) || (3'd6/*MS*/==-4'd7+xpc10nz) || (3'd6/*MS*/==-4'd6+xpc10nz) || (3'd6/*MS*/==-4'd5+xpc10nz) || (3'd6/*MS*/==
              -4'd4+xpc10nz) || (3'd6/*MS*/==-3'd3+xpc10nz) || (3'd6/*MS*/==-3'd2+xpc10nz) || (3'd6/*MS*/==-2'd1+xpc10nz) || (xpc10nz
              ==3'd6/*US*/)) && !xpc10_clear && !xpc10_stall;

               xpc10_trk5 <= ((3'd5/*MS*/==-11'd609+xpc10nz) || (3'd5/*MS*/==-11'd599+xpc10nz) || (3'd5/*MS*/==-11'd588+xpc10nz) || (3'd5
              /*MS*/==-11'd576+xpc10nz) || (3'd5/*MS*/==-11'd571+xpc10nz) || (3'd5/*MS*/==-11'd565+xpc10nz) || (3'd5/*MS*/==-11'd558+
              xpc10nz) || (3'd5/*MS*/==-11'd550+xpc10nz) || (3'd5/*MS*/==-11'd549+xpc10nz) || (3'd5/*MS*/==-11'd547+xpc10nz) || (3'd5
              /*MS*/==-11'd544+xpc10nz) || (3'd5/*MS*/==-11'd540+xpc10nz) || (3'd5/*MS*/==-11'd539+xpc10nz) || (3'd5/*MS*/==-11'd537+
              xpc10nz) || (3'd5/*MS*/==-11'd534+xpc10nz) || (3'd5/*MS*/==-11'd532+xpc10nz) || (3'd5/*MS*/==-11'd528+xpc10nz) || (3'd5
              /*MS*/==-10'd503+xpc10nz) || (3'd5/*MS*/==-10'd502+xpc10nz) || (3'd5/*MS*/==-10'd472+xpc10nz) || (3'd5/*MS*/==-10'd407+
              xpc10nz) || (3'd5/*MS*/==-10'd342+xpc10nz) || (3'd5/*MS*/==-10'd341+xpc10nz) || (3'd5/*MS*/==-10'd340+xpc10nz) || (3'd5
              /*MS*/==-10'd338+xpc10nz) || (3'd5/*MS*/==-10'd335+xpc10nz) || (3'd5/*MS*/==-10'd334+xpc10nz) || (3'd5/*MS*/==-10'd330+
              xpc10nz) || (3'd5/*MS*/==-10'd329+xpc10nz) || (3'd5/*MS*/==-10'd327+xpc10nz) || (3'd5/*MS*/==-10'd324+xpc10nz) || (3'd5
              /*MS*/==-10'd323+xpc10nz) || (3'd5/*MS*/==-10'd322+xpc10nz) || (3'd5/*MS*/==-10'd321+xpc10nz) || (3'd5/*MS*/==-10'd320+
              xpc10nz) || (3'd5/*MS*/==-10'd319+xpc10nz) || (3'd5/*MS*/==-10'd318+xpc10nz) || (3'd5/*MS*/==-10'd314+xpc10nz) || (3'd5
              /*MS*/==-10'd289+xpc10nz) || (3'd5/*MS*/==-10'd287+xpc10nz) || (3'd5/*MS*/==-10'd285+xpc10nz) || (3'd5/*MS*/==-10'd284+
              xpc10nz) || (3'd5/*MS*/==-10'd259+xpc10nz) || (3'd5/*MS*/==-10'd258+xpc10nz) || (3'd5/*MS*/==-10'd257+xpc10nz) || (3'd5
              /*MS*/==-9'd255+xpc10nz) || (3'd5/*MS*/==-9'd254+xpc10nz) || (3'd5/*MS*/==-9'd253+xpc10nz) || (3'd5/*MS*/==-9'd252+xpc10nz
              ) || (3'd5/*MS*/==-9'd251+xpc10nz) || (3'd5/*MS*/==-9'd250+xpc10nz) || (3'd5/*MS*/==-9'd249+xpc10nz) || (3'd5/*MS*/==-9'd248
              +xpc10nz) || (3'd5/*MS*/==-9'd247+xpc10nz) || (3'd5/*MS*/==-9'd246+xpc10nz) || (3'd5/*MS*/==-9'd245+xpc10nz) || (3'd5/*MS*/==
              -9'd244+xpc10nz) || (3'd5/*MS*/==-9'd242+xpc10nz) || (3'd5/*MS*/==-9'd241+xpc10nz) || (3'd5/*MS*/==-9'd239+xpc10nz) || 
              (3'd5/*MS*/==-9'd238+xpc10nz) || (3'd5/*MS*/==-9'd236+xpc10nz) || (3'd5/*MS*/==-9'd171+xpc10nz) || (3'd5/*MS*/==-8'd106
              +xpc10nz) || (3'd5/*MS*/==-8'd105+xpc10nz) || (3'd5/*MS*/==-8'd104+xpc10nz) || (3'd5/*MS*/==-8'd103+xpc10nz) || (3'd5/*MS*/==
              -8'd102+xpc10nz) || (3'd5/*MS*/==-8'd101+xpc10nz) || (3'd5/*MS*/==-8'd100+xpc10nz) || (3'd5/*MS*/==-8'd99+xpc10nz) || (3'd5
              /*MS*/==-8'd98+xpc10nz) || (3'd5/*MS*/==-8'd97+xpc10nz) || (3'd5/*MS*/==-8'd96+xpc10nz) || (3'd5/*MS*/==-8'd95+xpc10nz) || 
              (3'd5/*MS*/==-8'd94+xpc10nz) || (3'd5/*MS*/==-8'd93+xpc10nz) || (3'd5/*MS*/==-8'd92+xpc10nz) || (3'd5/*MS*/==-8'd91+xpc10nz
              ) || (3'd5/*MS*/==-8'd90+xpc10nz) || (3'd5/*MS*/==-8'd89+xpc10nz) || (3'd5/*MS*/==-8'd88+xpc10nz) || (3'd5/*MS*/==-8'd87
              +xpc10nz) || (3'd5/*MS*/==-8'd86+xpc10nz) || (3'd5/*MS*/==-8'd85+xpc10nz) || (3'd5/*MS*/==-8'd84+xpc10nz) || (3'd5/*MS*/==
              -8'd83+xpc10nz) || (3'd5/*MS*/==-8'd82+xpc10nz) || (3'd5/*MS*/==-8'd65+xpc10nz) || (3'd5/*MS*/==-8'd64+xpc10nz) || (3'd5
              /*MS*/==-7'd59+xpc10nz) || (3'd5/*MS*/==-7'd50+xpc10nz) || (3'd5/*MS*/==-7'd37+xpc10nz) || (3'd5/*MS*/==-6'd20+xpc10nz) || 
              (3'd5/*MS*/==-6'd19+xpc10nz) || (3'd5/*MS*/==-6'd18+xpc10nz) || (3'd5/*MS*/==-6'd17+xpc10nz) || (3'd5/*MS*/==-6'd16+xpc10nz
              ) || (3'd5/*MS*/==-5'd15+xpc10nz) || (3'd5/*MS*/==-5'd14+xpc10nz) || (3'd5/*MS*/==-5'd13+xpc10nz) || (3'd5/*MS*/==-5'd12
              +xpc10nz) || (3'd5/*MS*/==-5'd11+xpc10nz) || (3'd5/*MS*/==-5'd10+xpc10nz) || (3'd5/*MS*/==-5'd9+xpc10nz) || (3'd5/*MS*/==
              -5'd8+xpc10nz) || (3'd5/*MS*/==-4'd7+xpc10nz) || (3'd5/*MS*/==-4'd6+xpc10nz) || (3'd5/*MS*/==-4'd5+xpc10nz) || (3'd5/*MS*/==
              -4'd4+xpc10nz) || (3'd5/*MS*/==-3'd3+xpc10nz) || (3'd5/*MS*/==-3'd2+xpc10nz) || (3'd5/*MS*/==-2'd1+xpc10nz) || (xpc10nz
              ==3'd5/*US*/)) && !xpc10_clear && !xpc10_stall;

               xpc10_trk4 <= ((3'd4/*MS*/==-11'd609+xpc10nz) || (3'd4/*MS*/==-11'd599+xpc10nz) || (3'd4/*MS*/==-11'd588+xpc10nz) || (3'd4
              /*MS*/==-11'd576+xpc10nz) || (3'd4/*MS*/==-11'd571+xpc10nz) || (3'd4/*MS*/==-11'd565+xpc10nz) || (3'd4/*MS*/==-11'd558+
              xpc10nz) || (3'd4/*MS*/==-11'd550+xpc10nz) || (3'd4/*MS*/==-11'd549+xpc10nz) || (3'd4/*MS*/==-11'd547+xpc10nz) || (3'd4
              /*MS*/==-11'd544+xpc10nz) || (3'd4/*MS*/==-11'd540+xpc10nz) || (3'd4/*MS*/==-11'd539+xpc10nz) || (3'd4/*MS*/==-11'd537+
              xpc10nz) || (3'd4/*MS*/==-11'd534+xpc10nz) || (3'd4/*MS*/==-11'd532+xpc10nz) || (3'd4/*MS*/==-11'd528+xpc10nz) || (3'd4
              /*MS*/==-10'd503+xpc10nz) || (3'd4/*MS*/==-10'd502+xpc10nz) || (3'd4/*MS*/==-10'd472+xpc10nz) || (3'd4/*MS*/==-10'd407+
              xpc10nz) || (3'd4/*MS*/==-10'd342+xpc10nz) || (3'd4/*MS*/==-10'd341+xpc10nz) || (3'd4/*MS*/==-10'd340+xpc10nz) || (3'd4
              /*MS*/==-10'd338+xpc10nz) || (3'd4/*MS*/==-10'd335+xpc10nz) || (3'd4/*MS*/==-10'd334+xpc10nz) || (3'd4/*MS*/==-10'd330+
              xpc10nz) || (3'd4/*MS*/==-10'd329+xpc10nz) || (3'd4/*MS*/==-10'd327+xpc10nz) || (3'd4/*MS*/==-10'd324+xpc10nz) || (3'd4
              /*MS*/==-10'd323+xpc10nz) || (3'd4/*MS*/==-10'd322+xpc10nz) || (3'd4/*MS*/==-10'd321+xpc10nz) || (3'd4/*MS*/==-10'd320+
              xpc10nz) || (3'd4/*MS*/==-10'd319+xpc10nz) || (3'd4/*MS*/==-10'd318+xpc10nz) || (3'd4/*MS*/==-10'd314+xpc10nz) || (3'd4
              /*MS*/==-10'd289+xpc10nz) || (3'd4/*MS*/==-10'd287+xpc10nz) || (3'd4/*MS*/==-10'd285+xpc10nz) || (3'd4/*MS*/==-10'd284+
              xpc10nz) || (3'd4/*MS*/==-10'd259+xpc10nz) || (3'd4/*MS*/==-10'd258+xpc10nz) || (3'd4/*MS*/==-10'd257+xpc10nz) || (3'd4
              /*MS*/==-9'd255+xpc10nz) || (3'd4/*MS*/==-9'd254+xpc10nz) || (3'd4/*MS*/==-9'd253+xpc10nz) || (3'd4/*MS*/==-9'd252+xpc10nz
              ) || (3'd4/*MS*/==-9'd251+xpc10nz) || (3'd4/*MS*/==-9'd250+xpc10nz) || (3'd4/*MS*/==-9'd249+xpc10nz) || (3'd4/*MS*/==-9'd248
              +xpc10nz) || (3'd4/*MS*/==-9'd247+xpc10nz) || (3'd4/*MS*/==-9'd246+xpc10nz) || (3'd4/*MS*/==-9'd245+xpc10nz) || (3'd4/*MS*/==
              -9'd244+xpc10nz) || (3'd4/*MS*/==-9'd242+xpc10nz) || (3'd4/*MS*/==-9'd241+xpc10nz) || (3'd4/*MS*/==-9'd239+xpc10nz) || 
              (3'd4/*MS*/==-9'd238+xpc10nz) || (3'd4/*MS*/==-9'd236+xpc10nz) || (3'd4/*MS*/==-9'd171+xpc10nz) || (3'd4/*MS*/==-8'd106
              +xpc10nz) || (3'd4/*MS*/==-8'd105+xpc10nz) || (3'd4/*MS*/==-8'd104+xpc10nz) || (3'd4/*MS*/==-8'd103+xpc10nz) || (3'd4/*MS*/==
              -8'd102+xpc10nz) || (3'd4/*MS*/==-8'd101+xpc10nz) || (3'd4/*MS*/==-8'd100+xpc10nz) || (3'd4/*MS*/==-8'd99+xpc10nz) || (3'd4
              /*MS*/==-8'd98+xpc10nz) || (3'd4/*MS*/==-8'd97+xpc10nz) || (3'd4/*MS*/==-8'd96+xpc10nz) || (3'd4/*MS*/==-8'd95+xpc10nz) || 
              (3'd4/*MS*/==-8'd94+xpc10nz) || (3'd4/*MS*/==-8'd93+xpc10nz) || (3'd4/*MS*/==-8'd92+xpc10nz) || (3'd4/*MS*/==-8'd91+xpc10nz
              ) || (3'd4/*MS*/==-8'd90+xpc10nz) || (3'd4/*MS*/==-8'd89+xpc10nz) || (3'd4/*MS*/==-8'd88+xpc10nz) || (3'd4/*MS*/==-8'd87
              +xpc10nz) || (3'd4/*MS*/==-8'd86+xpc10nz) || (3'd4/*MS*/==-8'd85+xpc10nz) || (3'd4/*MS*/==-8'd84+xpc10nz) || (3'd4/*MS*/==
              -8'd83+xpc10nz) || (3'd4/*MS*/==-8'd82+xpc10nz) || (3'd4/*MS*/==-8'd65+xpc10nz) || (3'd4/*MS*/==-8'd64+xpc10nz) || (3'd4
              /*MS*/==-7'd59+xpc10nz) || (3'd4/*MS*/==-7'd50+xpc10nz) || (3'd4/*MS*/==-7'd37+xpc10nz) || (3'd4/*MS*/==-6'd20+xpc10nz) || 
              (3'd4/*MS*/==-6'd19+xpc10nz) || (3'd4/*MS*/==-6'd18+xpc10nz) || (3'd4/*MS*/==-6'd17+xpc10nz) || (3'd4/*MS*/==-6'd16+xpc10nz
              ) || (3'd4/*MS*/==-5'd15+xpc10nz) || (3'd4/*MS*/==-5'd14+xpc10nz) || (3'd4/*MS*/==-5'd13+xpc10nz) || (3'd4/*MS*/==-5'd12
              +xpc10nz) || (3'd4/*MS*/==-5'd11+xpc10nz) || (3'd4/*MS*/==-5'd10+xpc10nz) || (3'd4/*MS*/==-5'd9+xpc10nz) || (3'd4/*MS*/==
              -5'd8+xpc10nz) || (3'd4/*MS*/==-4'd7+xpc10nz) || (3'd4/*MS*/==-4'd6+xpc10nz) || (3'd4/*MS*/==-4'd5+xpc10nz) || (3'd4/*MS*/==
              -4'd4+xpc10nz) || (3'd4/*MS*/==-3'd3+xpc10nz) || (3'd4/*MS*/==-3'd2+xpc10nz) || (3'd4/*MS*/==-2'd1+xpc10nz) || (xpc10nz
              ==3'd4/*US*/)) && !xpc10_clear && !xpc10_stall;

               xpc10_trk3 <= ((2'd3/*MS*/==-11'd609+xpc10nz) || (2'd3/*MS*/==-11'd599+xpc10nz) || (2'd3/*MS*/==-11'd588+xpc10nz) || (2'd3
              /*MS*/==-11'd576+xpc10nz) || (2'd3/*MS*/==-11'd571+xpc10nz) || (2'd3/*MS*/==-11'd565+xpc10nz) || (2'd3/*MS*/==-11'd558+
              xpc10nz) || (2'd3/*MS*/==-11'd550+xpc10nz) || (2'd3/*MS*/==-11'd549+xpc10nz) || (2'd3/*MS*/==-11'd547+xpc10nz) || (2'd3
              /*MS*/==-11'd544+xpc10nz) || (2'd3/*MS*/==-11'd540+xpc10nz) || (2'd3/*MS*/==-11'd539+xpc10nz) || (2'd3/*MS*/==-11'd537+
              xpc10nz) || (2'd3/*MS*/==-11'd534+xpc10nz) || (2'd3/*MS*/==-11'd532+xpc10nz) || (2'd3/*MS*/==-11'd528+xpc10nz) || (2'd3
              /*MS*/==-10'd503+xpc10nz) || (2'd3/*MS*/==-10'd502+xpc10nz) || (2'd3/*MS*/==-10'd472+xpc10nz) || (2'd3/*MS*/==-10'd407+
              xpc10nz) || (2'd3/*MS*/==-10'd342+xpc10nz) || (2'd3/*MS*/==-10'd341+xpc10nz) || (2'd3/*MS*/==-10'd340+xpc10nz) || (2'd3
              /*MS*/==-10'd338+xpc10nz) || (2'd3/*MS*/==-10'd335+xpc10nz) || (2'd3/*MS*/==-10'd334+xpc10nz) || (2'd3/*MS*/==-10'd330+
              xpc10nz) || (2'd3/*MS*/==-10'd329+xpc10nz) || (2'd3/*MS*/==-10'd327+xpc10nz) || (2'd3/*MS*/==-10'd324+xpc10nz) || (2'd3
              /*MS*/==-10'd323+xpc10nz) || (2'd3/*MS*/==-10'd322+xpc10nz) || (2'd3/*MS*/==-10'd321+xpc10nz) || (2'd3/*MS*/==-10'd320+
              xpc10nz) || (2'd3/*MS*/==-10'd319+xpc10nz) || (2'd3/*MS*/==-10'd318+xpc10nz) || (2'd3/*MS*/==-10'd314+xpc10nz) || (2'd3
              /*MS*/==-10'd289+xpc10nz) || (2'd3/*MS*/==-10'd287+xpc10nz) || (2'd3/*MS*/==-10'd285+xpc10nz) || (2'd3/*MS*/==-10'd284+
              xpc10nz) || (2'd3/*MS*/==-10'd259+xpc10nz) || (2'd3/*MS*/==-10'd258+xpc10nz) || (2'd3/*MS*/==-10'd257+xpc10nz) || (2'd3
              /*MS*/==-9'd255+xpc10nz) || (2'd3/*MS*/==-9'd254+xpc10nz) || (2'd3/*MS*/==-9'd253+xpc10nz) || (2'd3/*MS*/==-9'd252+xpc10nz
              ) || (2'd3/*MS*/==-9'd251+xpc10nz) || (2'd3/*MS*/==-9'd250+xpc10nz) || (2'd3/*MS*/==-9'd249+xpc10nz) || (2'd3/*MS*/==-9'd248
              +xpc10nz) || (2'd3/*MS*/==-9'd247+xpc10nz) || (2'd3/*MS*/==-9'd246+xpc10nz) || (2'd3/*MS*/==-9'd245+xpc10nz) || (2'd3/*MS*/==
              -9'd244+xpc10nz) || (2'd3/*MS*/==-9'd242+xpc10nz) || (2'd3/*MS*/==-9'd241+xpc10nz) || (2'd3/*MS*/==-9'd239+xpc10nz) || 
              (2'd3/*MS*/==-9'd238+xpc10nz) || (2'd3/*MS*/==-9'd236+xpc10nz) || (2'd3/*MS*/==-9'd171+xpc10nz) || (2'd3/*MS*/==-8'd106
              +xpc10nz) || (2'd3/*MS*/==-8'd105+xpc10nz) || (2'd3/*MS*/==-8'd104+xpc10nz) || (2'd3/*MS*/==-8'd103+xpc10nz) || (2'd3/*MS*/==
              -8'd102+xpc10nz) || (2'd3/*MS*/==-8'd101+xpc10nz) || (2'd3/*MS*/==-8'd100+xpc10nz) || (2'd3/*MS*/==-8'd99+xpc10nz) || (2'd3
              /*MS*/==-8'd98+xpc10nz) || (2'd3/*MS*/==-8'd97+xpc10nz) || (2'd3/*MS*/==-8'd96+xpc10nz) || (2'd3/*MS*/==-8'd95+xpc10nz) || 
              (2'd3/*MS*/==-8'd94+xpc10nz) || (2'd3/*MS*/==-8'd93+xpc10nz) || (2'd3/*MS*/==-8'd92+xpc10nz) || (2'd3/*MS*/==-8'd91+xpc10nz
              ) || (2'd3/*MS*/==-8'd90+xpc10nz) || (2'd3/*MS*/==-8'd89+xpc10nz) || (2'd3/*MS*/==-8'd88+xpc10nz) || (2'd3/*MS*/==-8'd87
              +xpc10nz) || (2'd3/*MS*/==-8'd86+xpc10nz) || (2'd3/*MS*/==-8'd85+xpc10nz) || (2'd3/*MS*/==-8'd84+xpc10nz) || (2'd3/*MS*/==
              -8'd83+xpc10nz) || (2'd3/*MS*/==-8'd82+xpc10nz) || (2'd3/*MS*/==-8'd65+xpc10nz) || (2'd3/*MS*/==-8'd64+xpc10nz) || (2'd3
              /*MS*/==-7'd59+xpc10nz) || (2'd3/*MS*/==-7'd50+xpc10nz) || (2'd3/*MS*/==-7'd37+xpc10nz) || (2'd3/*MS*/==-6'd20+xpc10nz) || 
              (2'd3/*MS*/==-6'd19+xpc10nz) || (2'd3/*MS*/==-6'd18+xpc10nz) || (2'd3/*MS*/==-6'd17+xpc10nz) || (2'd3/*MS*/==-6'd16+xpc10nz
              ) || (2'd3/*MS*/==-5'd15+xpc10nz) || (2'd3/*MS*/==-5'd14+xpc10nz) || (2'd3/*MS*/==-5'd13+xpc10nz) || (2'd3/*MS*/==-5'd12
              +xpc10nz) || (2'd3/*MS*/==-5'd11+xpc10nz) || (2'd3/*MS*/==-5'd10+xpc10nz) || (2'd3/*MS*/==-5'd9+xpc10nz) || (2'd3/*MS*/==
              -5'd8+xpc10nz) || (2'd3/*MS*/==-4'd7+xpc10nz) || (2'd3/*MS*/==-4'd6+xpc10nz) || (2'd3/*MS*/==-4'd5+xpc10nz) || (2'd3/*MS*/==
              -4'd4+xpc10nz) || (2'd3/*MS*/==-3'd3+xpc10nz) || (2'd3/*MS*/==-3'd2+xpc10nz) || (2'd3/*MS*/==-2'd1+xpc10nz) || (xpc10nz
              ==2'd3/*US*/)) && !xpc10_clear && !xpc10_stall;

               xpc10_trk2 <= ((2'd2/*MS*/==-11'd609+xpc10nz) || (2'd2/*MS*/==-11'd599+xpc10nz) || (2'd2/*MS*/==-11'd588+xpc10nz) || (2'd2
              /*MS*/==-11'd576+xpc10nz) || (2'd2/*MS*/==-11'd571+xpc10nz) || (2'd2/*MS*/==-11'd565+xpc10nz) || (2'd2/*MS*/==-11'd558+
              xpc10nz) || (2'd2/*MS*/==-11'd550+xpc10nz) || (2'd2/*MS*/==-11'd549+xpc10nz) || (2'd2/*MS*/==-11'd547+xpc10nz) || (2'd2
              /*MS*/==-11'd544+xpc10nz) || (2'd2/*MS*/==-11'd540+xpc10nz) || (2'd2/*MS*/==-11'd539+xpc10nz) || (2'd2/*MS*/==-11'd537+
              xpc10nz) || (2'd2/*MS*/==-11'd534+xpc10nz) || (2'd2/*MS*/==-11'd532+xpc10nz) || (2'd2/*MS*/==-11'd528+xpc10nz) || (2'd2
              /*MS*/==-10'd503+xpc10nz) || (2'd2/*MS*/==-10'd502+xpc10nz) || (2'd2/*MS*/==-10'd472+xpc10nz) || (2'd2/*MS*/==-10'd407+
              xpc10nz) || (2'd2/*MS*/==-10'd342+xpc10nz) || (2'd2/*MS*/==-10'd341+xpc10nz) || (2'd2/*MS*/==-10'd340+xpc10nz) || (2'd2
              /*MS*/==-10'd338+xpc10nz) || (2'd2/*MS*/==-10'd335+xpc10nz) || (2'd2/*MS*/==-10'd334+xpc10nz) || (2'd2/*MS*/==-10'd330+
              xpc10nz) || (2'd2/*MS*/==-10'd329+xpc10nz) || (2'd2/*MS*/==-10'd327+xpc10nz) || (2'd2/*MS*/==-10'd324+xpc10nz) || (2'd2
              /*MS*/==-10'd323+xpc10nz) || (2'd2/*MS*/==-10'd322+xpc10nz) || (2'd2/*MS*/==-10'd321+xpc10nz) || (2'd2/*MS*/==-10'd320+
              xpc10nz) || (2'd2/*MS*/==-10'd319+xpc10nz) || (2'd2/*MS*/==-10'd318+xpc10nz) || (2'd2/*MS*/==-10'd314+xpc10nz) || (2'd2
              /*MS*/==-10'd289+xpc10nz) || (2'd2/*MS*/==-10'd287+xpc10nz) || (2'd2/*MS*/==-10'd285+xpc10nz) || (2'd2/*MS*/==-10'd284+
              xpc10nz) || (2'd2/*MS*/==-10'd259+xpc10nz) || (2'd2/*MS*/==-10'd258+xpc10nz) || (2'd2/*MS*/==-10'd257+xpc10nz) || (2'd2
              /*MS*/==-9'd255+xpc10nz) || (2'd2/*MS*/==-9'd254+xpc10nz) || (2'd2/*MS*/==-9'd253+xpc10nz) || (2'd2/*MS*/==-9'd252+xpc10nz
              ) || (2'd2/*MS*/==-9'd251+xpc10nz) || (2'd2/*MS*/==-9'd250+xpc10nz) || (2'd2/*MS*/==-9'd249+xpc10nz) || (2'd2/*MS*/==-9'd248
              +xpc10nz) || (2'd2/*MS*/==-9'd247+xpc10nz) || (2'd2/*MS*/==-9'd246+xpc10nz) || (2'd2/*MS*/==-9'd245+xpc10nz) || (2'd2/*MS*/==
              -9'd244+xpc10nz) || (2'd2/*MS*/==-9'd242+xpc10nz) || (2'd2/*MS*/==-9'd241+xpc10nz) || (2'd2/*MS*/==-9'd239+xpc10nz) || 
              (2'd2/*MS*/==-9'd238+xpc10nz) || (2'd2/*MS*/==-9'd236+xpc10nz) || (2'd2/*MS*/==-9'd171+xpc10nz) || (2'd2/*MS*/==-8'd106
              +xpc10nz) || (2'd2/*MS*/==-8'd105+xpc10nz) || (2'd2/*MS*/==-8'd104+xpc10nz) || (2'd2/*MS*/==-8'd103+xpc10nz) || (2'd2/*MS*/==
              -8'd102+xpc10nz) || (2'd2/*MS*/==-8'd101+xpc10nz) || (2'd2/*MS*/==-8'd100+xpc10nz) || (2'd2/*MS*/==-8'd99+xpc10nz) || (2'd2
              /*MS*/==-8'd98+xpc10nz) || (2'd2/*MS*/==-8'd97+xpc10nz) || (2'd2/*MS*/==-8'd96+xpc10nz) || (2'd2/*MS*/==-8'd95+xpc10nz) || 
              (2'd2/*MS*/==-8'd94+xpc10nz) || (2'd2/*MS*/==-8'd93+xpc10nz) || (2'd2/*MS*/==-8'd92+xpc10nz) || (2'd2/*MS*/==-8'd91+xpc10nz
              ) || (2'd2/*MS*/==-8'd90+xpc10nz) || (2'd2/*MS*/==-8'd89+xpc10nz) || (2'd2/*MS*/==-8'd88+xpc10nz) || (2'd2/*MS*/==-8'd87
              +xpc10nz) || (2'd2/*MS*/==-8'd86+xpc10nz) || (2'd2/*MS*/==-8'd85+xpc10nz) || (2'd2/*MS*/==-8'd84+xpc10nz) || (2'd2/*MS*/==
              -8'd83+xpc10nz) || (2'd2/*MS*/==-8'd82+xpc10nz) || (2'd2/*MS*/==-8'd65+xpc10nz) || (2'd2/*MS*/==-8'd64+xpc10nz) || (2'd2
              /*MS*/==-7'd59+xpc10nz) || (2'd2/*MS*/==-7'd50+xpc10nz) || (2'd2/*MS*/==-7'd37+xpc10nz) || (2'd2/*MS*/==-6'd20+xpc10nz) || 
              (2'd2/*MS*/==-6'd19+xpc10nz) || (2'd2/*MS*/==-6'd18+xpc10nz) || (2'd2/*MS*/==-6'd17+xpc10nz) || (2'd2/*MS*/==-6'd16+xpc10nz
              ) || (2'd2/*MS*/==-5'd15+xpc10nz) || (2'd2/*MS*/==-5'd14+xpc10nz) || (2'd2/*MS*/==-5'd13+xpc10nz) || (2'd2/*MS*/==-5'd12
              +xpc10nz) || (2'd2/*MS*/==-5'd11+xpc10nz) || (2'd2/*MS*/==-5'd10+xpc10nz) || (2'd2/*MS*/==-5'd9+xpc10nz) || (2'd2/*MS*/==
              -5'd8+xpc10nz) || (2'd2/*MS*/==-4'd7+xpc10nz) || (2'd2/*MS*/==-4'd6+xpc10nz) || (2'd2/*MS*/==-4'd5+xpc10nz) || (2'd2/*MS*/==
              -4'd4+xpc10nz) || (2'd2/*MS*/==-3'd3+xpc10nz) || (2'd2/*MS*/==-3'd2+xpc10nz) || (2'd2/*MS*/==-2'd1+xpc10nz) || (xpc10nz
              ==2'd2/*US*/)) && !xpc10_clear && !xpc10_stall;

               xpc10_trk1 <= ((1'd1/*MS*/==-11'd609+xpc10nz) || (1'd1/*MS*/==-11'd599+xpc10nz) || (1'd1/*MS*/==-11'd588+xpc10nz) || (1'd1
              /*MS*/==-11'd576+xpc10nz) || (1'd1/*MS*/==-11'd571+xpc10nz) || (1'd1/*MS*/==-11'd565+xpc10nz) || (1'd1/*MS*/==-11'd558+
              xpc10nz) || (1'd1/*MS*/==-11'd550+xpc10nz) || (1'd1/*MS*/==-11'd549+xpc10nz) || (1'd1/*MS*/==-11'd547+xpc10nz) || (1'd1
              /*MS*/==-11'd544+xpc10nz) || (1'd1/*MS*/==-11'd540+xpc10nz) || (1'd1/*MS*/==-11'd539+xpc10nz) || (1'd1/*MS*/==-11'd537+
              xpc10nz) || (1'd1/*MS*/==-11'd534+xpc10nz) || (1'd1/*MS*/==-11'd532+xpc10nz) || (1'd1/*MS*/==-11'd528+xpc10nz) || (1'd1
              /*MS*/==-10'd503+xpc10nz) || (1'd1/*MS*/==-10'd502+xpc10nz) || (1'd1/*MS*/==-10'd472+xpc10nz) || (1'd1/*MS*/==-10'd407+
              xpc10nz) || (1'd1/*MS*/==-10'd342+xpc10nz) || (1'd1/*MS*/==-10'd341+xpc10nz) || (1'd1/*MS*/==-10'd340+xpc10nz) || (1'd1
              /*MS*/==-10'd338+xpc10nz) || (1'd1/*MS*/==-10'd335+xpc10nz) || (1'd1/*MS*/==-10'd334+xpc10nz) || (1'd1/*MS*/==-10'd330+
              xpc10nz) || (1'd1/*MS*/==-10'd329+xpc10nz) || (1'd1/*MS*/==-10'd327+xpc10nz) || (1'd1/*MS*/==-10'd324+xpc10nz) || (1'd1
              /*MS*/==-10'd323+xpc10nz) || (1'd1/*MS*/==-10'd322+xpc10nz) || (1'd1/*MS*/==-10'd321+xpc10nz) || (1'd1/*MS*/==-10'd320+
              xpc10nz) || (1'd1/*MS*/==-10'd319+xpc10nz) || (1'd1/*MS*/==-10'd318+xpc10nz) || (1'd1/*MS*/==-10'd314+xpc10nz) || (1'd1
              /*MS*/==-10'd289+xpc10nz) || (1'd1/*MS*/==-10'd287+xpc10nz) || (1'd1/*MS*/==-10'd285+xpc10nz) || (1'd1/*MS*/==-10'd284+
              xpc10nz) || (1'd1/*MS*/==-10'd259+xpc10nz) || (1'd1/*MS*/==-10'd258+xpc10nz) || (1'd1/*MS*/==-10'd257+xpc10nz) || (1'd1
              /*MS*/==-9'd255+xpc10nz) || (1'd1/*MS*/==-9'd254+xpc10nz) || (1'd1/*MS*/==-9'd253+xpc10nz) || (1'd1/*MS*/==-9'd252+xpc10nz
              ) || (1'd1/*MS*/==-9'd251+xpc10nz) || (1'd1/*MS*/==-9'd250+xpc10nz) || (1'd1/*MS*/==-9'd249+xpc10nz) || (1'd1/*MS*/==-9'd248
              +xpc10nz) || (1'd1/*MS*/==-9'd247+xpc10nz) || (1'd1/*MS*/==-9'd246+xpc10nz) || (1'd1/*MS*/==-9'd245+xpc10nz) || (1'd1/*MS*/==
              -9'd244+xpc10nz) || (1'd1/*MS*/==-9'd242+xpc10nz) || (1'd1/*MS*/==-9'd241+xpc10nz) || (1'd1/*MS*/==-9'd239+xpc10nz) || 
              (1'd1/*MS*/==-9'd238+xpc10nz) || (1'd1/*MS*/==-9'd236+xpc10nz) || (1'd1/*MS*/==-9'd171+xpc10nz) || (1'd1/*MS*/==-8'd106
              +xpc10nz) || (1'd1/*MS*/==-8'd105+xpc10nz) || (1'd1/*MS*/==-8'd104+xpc10nz) || (1'd1/*MS*/==-8'd103+xpc10nz) || (1'd1/*MS*/==
              -8'd102+xpc10nz) || (1'd1/*MS*/==-8'd101+xpc10nz) || (1'd1/*MS*/==-8'd100+xpc10nz) || (1'd1/*MS*/==-8'd99+xpc10nz) || (1'd1
              /*MS*/==-8'd98+xpc10nz) || (1'd1/*MS*/==-8'd97+xpc10nz) || (1'd1/*MS*/==-8'd96+xpc10nz) || (1'd1/*MS*/==-8'd95+xpc10nz) || 
              (1'd1/*MS*/==-8'd94+xpc10nz) || (1'd1/*MS*/==-8'd93+xpc10nz) || (1'd1/*MS*/==-8'd92+xpc10nz) || (1'd1/*MS*/==-8'd91+xpc10nz
              ) || (1'd1/*MS*/==-8'd90+xpc10nz) || (1'd1/*MS*/==-8'd89+xpc10nz) || (1'd1/*MS*/==-8'd88+xpc10nz) || (1'd1/*MS*/==-8'd87
              +xpc10nz) || (1'd1/*MS*/==-8'd86+xpc10nz) || (1'd1/*MS*/==-8'd85+xpc10nz) || (1'd1/*MS*/==-8'd84+xpc10nz) || (1'd1/*MS*/==
              -8'd83+xpc10nz) || (1'd1/*MS*/==-8'd82+xpc10nz) || (1'd1/*MS*/==-8'd65+xpc10nz) || (1'd1/*MS*/==-8'd64+xpc10nz) || (1'd1
              /*MS*/==-7'd59+xpc10nz) || (1'd1/*MS*/==-7'd50+xpc10nz) || (1'd1/*MS*/==-7'd37+xpc10nz) || (1'd1/*MS*/==-6'd20+xpc10nz) || 
              (1'd1/*MS*/==-6'd19+xpc10nz) || (1'd1/*MS*/==-6'd18+xpc10nz) || (1'd1/*MS*/==-6'd17+xpc10nz) || (1'd1/*MS*/==-6'd16+xpc10nz
              ) || (1'd1/*MS*/==-5'd15+xpc10nz) || (1'd1/*MS*/==-5'd14+xpc10nz) || (1'd1/*MS*/==-5'd13+xpc10nz) || (1'd1/*MS*/==-5'd12
              +xpc10nz) || (1'd1/*MS*/==-5'd11+xpc10nz) || (1'd1/*MS*/==-5'd10+xpc10nz) || (1'd1/*MS*/==-5'd9+xpc10nz) || (1'd1/*MS*/==
              -5'd8+xpc10nz) || (1'd1/*MS*/==-4'd7+xpc10nz) || (1'd1/*MS*/==-4'd6+xpc10nz) || (1'd1/*MS*/==-4'd5+xpc10nz) || (1'd1/*MS*/==
              -4'd4+xpc10nz) || (1'd1/*MS*/==-3'd3+xpc10nz) || (1'd1/*MS*/==-3'd2+xpc10nz) || (1'd1/*MS*/==-2'd1+xpc10nz) || (xpc10nz
              ==1'd1/*US*/)) && !xpc10_clear && !xpc10_stall;

               xpc10_trk0 <= ((0/*MS*/==-11'd609+xpc10nz) || (0/*MS*/==-11'd599+xpc10nz) || (0/*MS*/==-11'd588+xpc10nz) || (0/*MS*/==
              -11'd576+xpc10nz) || (0/*MS*/==-11'd571+xpc10nz) || (0/*MS*/==-11'd565+xpc10nz) || (0/*MS*/==-11'd558+xpc10nz) || (0/*MS*/==
              -11'd550+xpc10nz) || (0/*MS*/==-11'd549+xpc10nz) || (0/*MS*/==-11'd547+xpc10nz) || (0/*MS*/==-11'd544+xpc10nz) || (0/*MS*/==
              -11'd540+xpc10nz) || (0/*MS*/==-11'd539+xpc10nz) || (0/*MS*/==-11'd537+xpc10nz) || (0/*MS*/==-11'd534+xpc10nz) || (0/*MS*/==
              -11'd532+xpc10nz) || (0/*MS*/==-11'd528+xpc10nz) || (0/*MS*/==-10'd503+xpc10nz) || (0/*MS*/==-10'd502+xpc10nz) || (0/*MS*/==
              -10'd472+xpc10nz) || (0/*MS*/==-10'd407+xpc10nz) || (0/*MS*/==-10'd342+xpc10nz) || (0/*MS*/==-10'd341+xpc10nz) || (0/*MS*/==
              -10'd340+xpc10nz) || (0/*MS*/==-10'd338+xpc10nz) || (0/*MS*/==-10'd335+xpc10nz) || (0/*MS*/==-10'd334+xpc10nz) || (0/*MS*/==
              -10'd330+xpc10nz) || (0/*MS*/==-10'd329+xpc10nz) || (0/*MS*/==-10'd327+xpc10nz) || (0/*MS*/==-10'd324+xpc10nz) || (0/*MS*/==
              -10'd323+xpc10nz) || (0/*MS*/==-10'd322+xpc10nz) || (0/*MS*/==-10'd321+xpc10nz) || (0/*MS*/==-10'd320+xpc10nz) || (0/*MS*/==
              -10'd319+xpc10nz) || (0/*MS*/==-10'd318+xpc10nz) || (0/*MS*/==-10'd314+xpc10nz) || (0/*MS*/==-10'd289+xpc10nz) || (0/*MS*/==
              -10'd287+xpc10nz) || (0/*MS*/==-10'd285+xpc10nz) || (0/*MS*/==-10'd284+xpc10nz) || (0/*MS*/==-10'd259+xpc10nz) || (0/*MS*/==
              -10'd258+xpc10nz) || (0/*MS*/==-10'd257+xpc10nz) || (0/*MS*/==-9'd255+xpc10nz) || (0/*MS*/==-9'd254+xpc10nz) || (0/*MS*/==
              -9'd253+xpc10nz) || (0/*MS*/==-9'd252+xpc10nz) || (0/*MS*/==-9'd251+xpc10nz) || (0/*MS*/==-9'd250+xpc10nz) || (0/*MS*/==
              -9'd249+xpc10nz) || (0/*MS*/==-9'd248+xpc10nz) || (0/*MS*/==-9'd247+xpc10nz) || (0/*MS*/==-9'd246+xpc10nz) || (0/*MS*/==
              -9'd245+xpc10nz) || (0/*MS*/==-9'd244+xpc10nz) || (0/*MS*/==-9'd242+xpc10nz) || (0/*MS*/==-9'd241+xpc10nz) || (0/*MS*/==
              -9'd239+xpc10nz) || (0/*MS*/==-9'd238+xpc10nz) || (0/*MS*/==-9'd236+xpc10nz) || (0/*MS*/==-9'd171+xpc10nz) || (0/*MS*/==
              -8'd106+xpc10nz) || (0/*MS*/==-8'd105+xpc10nz) || (0/*MS*/==-8'd104+xpc10nz) || (0/*MS*/==-8'd103+xpc10nz) || (0/*MS*/==
              -8'd102+xpc10nz) || (0/*MS*/==-8'd101+xpc10nz) || (0/*MS*/==-8'd100+xpc10nz) || (0/*MS*/==-8'd99+xpc10nz) || (0/*MS*/==
              -8'd98+xpc10nz) || (0/*MS*/==-8'd97+xpc10nz) || (0/*MS*/==-8'd96+xpc10nz) || (0/*MS*/==-8'd95+xpc10nz) || (0/*MS*/==-8'd94
              +xpc10nz) || (0/*MS*/==-8'd93+xpc10nz) || (0/*MS*/==-8'd92+xpc10nz) || (0/*MS*/==-8'd91+xpc10nz) || (0/*MS*/==-8'd90+xpc10nz
              ) || (0/*MS*/==-8'd89+xpc10nz) || (0/*MS*/==-8'd88+xpc10nz) || (0/*MS*/==-8'd87+xpc10nz) || (0/*MS*/==-8'd86+xpc10nz) || 
              (0/*MS*/==-8'd85+xpc10nz) || (0/*MS*/==-8'd84+xpc10nz) || (0/*MS*/==-8'd83+xpc10nz) || (0/*MS*/==-8'd82+xpc10nz) || (0/*MS*/==
              -8'd65+xpc10nz) || (0/*MS*/==-8'd64+xpc10nz) || (0/*MS*/==-7'd59+xpc10nz) || (0/*MS*/==-7'd50+xpc10nz) || (0/*MS*/==-7'd37
              +xpc10nz) || (0/*MS*/==-6'd20+xpc10nz) || (0/*MS*/==-6'd19+xpc10nz) || (0/*MS*/==-6'd18+xpc10nz) || (0/*MS*/==-6'd17+xpc10nz
              ) || (0/*MS*/==-6'd16+xpc10nz) || (0/*MS*/==-5'd15+xpc10nz) || (0/*MS*/==-5'd14+xpc10nz) || (0/*MS*/==-5'd13+xpc10nz) || 
              (0/*MS*/==-5'd12+xpc10nz) || (0/*MS*/==-5'd11+xpc10nz) || (0/*MS*/==-5'd10+xpc10nz) || (0/*MS*/==-5'd9+xpc10nz) || (0/*MS*/==
              -5'd8+xpc10nz) || (0/*MS*/==-4'd7+xpc10nz) || (0/*MS*/==-4'd6+xpc10nz) || (0/*MS*/==-4'd5+xpc10nz) || (0/*MS*/==-4'd4+xpc10nz
              ) || (0/*MS*/==-3'd3+xpc10nz) || (0/*MS*/==-3'd2+xpc10nz) || (0/*MS*/==-2'd1+xpc10nz) || (xpc10nz==0/*US*/)) && !xpc10_clear
               && !xpc10_stall;

              if ((xpc10nz==0/*US*/))  xpc10nz <= 1'd1/*xpc10nz*/;
                  if ((xpc10nz==2'd2/*US*/))  xpc10nz <= 2'd3/*US*/;
                  if ((xpc10nz==2'd3/*US*/))  xpc10nz <= 3'd4/*xpc10nz*/;
                  if ((xpc10nz==3'd6/*US*/))  xpc10nz <= 3'd7/*xpc10nz*/;
                  if ((xpc10nz==4'd9/*US*/))  xpc10nz <= 4'd10/*xpc10nz*/;
                  if ((xpc10nz==4'd11/*US*/))  xpc10nz <= 4'd12/*xpc10nz*/;
                  if ((xpc10nz==4'd14/*US*/))  xpc10nz <= 4'd15/*xpc10nz*/;
                  if ((xpc10nz==5'd17/*US*/))  xpc10nz <= 5'd18/*US*/;
                  if ((xpc10nz==5'd18/*US*/))  xpc10nz <= 5'd19/*xpc10nz*/;
                  if ((xpc10nz==5'd21/*US*/))  xpc10nz <= 6'd37/*xpc10nz*/;
                  if ((xpc10nz==5'd22/*US*/))  xpc10nz <= 6'd37/*xpc10nz*/;
                  if ((xpc10nz==5'd23/*US*/))  xpc10nz <= 6'd37/*xpc10nz*/;
                  if ((xpc10nz==5'd24/*US*/))  xpc10nz <= 6'd37/*xpc10nz*/;
                  if ((xpc10nz==5'd25/*US*/))  xpc10nz <= 10'd576/*xpc10nz*/;
                  if ((xpc10nz==5'd26/*US*/))  xpc10nz <= 10'd588/*xpc10nz*/;
                  if ((xpc10nz==5'd27/*US*/))  xpc10nz <= 10'd599/*xpc10nz*/;
                  if ((xpc10nz==5'd28/*US*/))  xpc10nz <= 10'd609/*xpc10nz*/;
                  if ((xpc10nz==5'd29/*US*/))  xpc10nz <= 10'd550/*xpc10nz*/;
                  if ((xpc10nz==5'd30/*US*/))  xpc10nz <= 10'd558/*xpc10nz*/;
                  if ((xpc10nz==5'd31/*US*/))  xpc10nz <= 10'd565/*xpc10nz*/;
                  if ((xpc10nz==6'd32/*US*/))  xpc10nz <= 10'd571/*xpc10nz*/;
                  if ((xpc10nz==6'd33/*US*/))  xpc10nz <= 10'd540/*xpc10nz*/;
                  if ((xpc10nz==6'd34/*US*/))  xpc10nz <= 10'd544/*xpc10nz*/;
                  if ((xpc10nz==6'd35/*US*/))  xpc10nz <= 10'd547/*xpc10nz*/;
                  if ((xpc10nz==6'd36/*US*/))  xpc10nz <= 10'd549/*xpc10nz*/;
                  if ((xpc10nz==6'd38/*US*/))  xpc10nz <= 6'd50/*xpc10nz*/;
                  if ((xpc10nz==6'd39/*US*/))  xpc10nz <= 6'd50/*xpc10nz*/;
                  if ((xpc10nz==6'd40/*US*/))  xpc10nz <= 6'd50/*xpc10nz*/;
                  if ((xpc10nz==6'd41/*US*/))  xpc10nz <= 6'd50/*xpc10nz*/;
                  if ((xpc10nz==6'd42/*US*/))  xpc10nz <= 10'd550/*xpc10nz*/;
                  if ((xpc10nz==6'd43/*US*/))  xpc10nz <= 10'd558/*xpc10nz*/;
                  if ((xpc10nz==6'd44/*US*/))  xpc10nz <= 10'd565/*xpc10nz*/;
                  if ((xpc10nz==6'd45/*US*/))  xpc10nz <= 10'd571/*xpc10nz*/;
                  if ((xpc10nz==6'd46/*US*/))  xpc10nz <= 10'd540/*xpc10nz*/;
                  if ((xpc10nz==6'd47/*US*/))  xpc10nz <= 10'd544/*xpc10nz*/;
                  if ((xpc10nz==6'd48/*US*/))  xpc10nz <= 10'd547/*xpc10nz*/;
                  if ((xpc10nz==6'd49/*US*/))  xpc10nz <= 10'd549/*xpc10nz*/;
                  if ((xpc10nz==6'd51/*US*/))  xpc10nz <= 6'd59/*xpc10nz*/;
                  if ((xpc10nz==6'd52/*US*/))  xpc10nz <= 6'd59/*xpc10nz*/;
                  if ((xpc10nz==6'd53/*US*/))  xpc10nz <= 6'd59/*xpc10nz*/;
                  if ((xpc10nz==6'd54/*US*/))  xpc10nz <= 6'd59/*xpc10nz*/;
                  if ((xpc10nz==6'd55/*US*/))  xpc10nz <= 10'd540/*xpc10nz*/;
                  if ((xpc10nz==6'd56/*US*/))  xpc10nz <= 10'd544/*xpc10nz*/;
                  if ((xpc10nz==6'd57/*US*/))  xpc10nz <= 10'd547/*xpc10nz*/;
                  if ((xpc10nz==6'd58/*US*/))  xpc10nz <= 10'd549/*xpc10nz*/;
                  if ((xpc10nz==6'd60/*US*/))  xpc10nz <= 7'd64/*xpc10nz*/;
                  if ((xpc10nz==6'd61/*US*/))  xpc10nz <= 7'd64/*xpc10nz*/;
                  if ((xpc10nz==6'd62/*US*/))  xpc10nz <= 7'd64/*xpc10nz*/;
                  if ((xpc10nz==6'd63/*US*/))  xpc10nz <= 7'd64/*xpc10nz*/;
                  if ((xpc10nz==7'd66/*US*/))  xpc10nz <= 10'd528/*xpc10nz*/;
                  if ((xpc10nz==7'd67/*US*/))  xpc10nz <= 10'd534/*xpc10nz*/;
                  if ((xpc10nz==7'd68/*US*/))  xpc10nz <= 10'd537/*xpc10nz*/;
                  if ((xpc10nz==7'd69/*US*/))  xpc10nz <= 10'd539/*xpc10nz*/;
                  if ((xpc10nz==7'd70/*US*/))  xpc10nz <= 10'd528/*xpc10nz*/;
                  if ((xpc10nz==7'd71/*US*/))  xpc10nz <= 10'd534/*xpc10nz*/;
                  if ((xpc10nz==7'd72/*US*/))  xpc10nz <= 10'd537/*xpc10nz*/;
                  if ((xpc10nz==7'd73/*US*/))  xpc10nz <= 10'd539/*xpc10nz*/;
                  if ((xpc10nz==7'd74/*US*/))  xpc10nz <= 10'd528/*xpc10nz*/;
                  if ((xpc10nz==7'd75/*US*/))  xpc10nz <= 10'd534/*xpc10nz*/;
                  if ((xpc10nz==7'd76/*US*/))  xpc10nz <= 10'd537/*xpc10nz*/;
                  if ((xpc10nz==7'd77/*US*/))  xpc10nz <= 10'd539/*xpc10nz*/;
                  if ((xpc10nz==7'd78/*US*/))  xpc10nz <= 10'd528/*xpc10nz*/;
                  if ((xpc10nz==7'd79/*US*/))  xpc10nz <= 10'd534/*xpc10nz*/;
                  if ((xpc10nz==7'd80/*US*/))  xpc10nz <= 10'd537/*xpc10nz*/;
                  if ((xpc10nz==7'd81/*US*/))  xpc10nz <= 10'd539/*xpc10nz*/;
                  if ((xpc10nz==7'd107/*US*/))  xpc10nz <= 7'd108/*xpc10nz*/;
                  if ((xpc10nz==7'd108/*US*/))  xpc10nz <= 7'd109/*xpc10nz*/;
                  if ((xpc10nz==7'd109/*US*/))  xpc10nz <= 7'd110/*xpc10nz*/;
                  if ((xpc10nz==7'd110/*US*/))  xpc10nz <= 7'd111/*xpc10nz*/;
                  if ((xpc10nz==7'd111/*US*/))  xpc10nz <= 7'd112/*xpc10nz*/;
                  if ((xpc10nz==7'd112/*US*/))  xpc10nz <= 7'd113/*xpc10nz*/;
                  if ((xpc10nz==7'd113/*US*/))  xpc10nz <= 7'd114/*xpc10nz*/;
                  if ((xpc10nz==7'd114/*US*/))  xpc10nz <= 7'd115/*xpc10nz*/;
                  if ((xpc10nz==7'd115/*US*/))  xpc10nz <= 7'd116/*xpc10nz*/;
                  if ((xpc10nz==7'd116/*US*/))  xpc10nz <= 7'd117/*xpc10nz*/;
                  if ((xpc10nz==7'd117/*US*/))  xpc10nz <= 7'd118/*xpc10nz*/;
                  if ((xpc10nz==7'd118/*US*/))  xpc10nz <= 7'd119/*xpc10nz*/;
                  if ((xpc10nz==7'd119/*US*/))  xpc10nz <= 7'd120/*xpc10nz*/;
                  if ((xpc10nz==7'd120/*US*/))  xpc10nz <= 7'd121/*xpc10nz*/;
                  if ((xpc10nz==7'd121/*US*/))  xpc10nz <= 7'd122/*xpc10nz*/;
                  if ((xpc10nz==7'd122/*US*/))  xpc10nz <= 7'd123/*xpc10nz*/;
                  if ((xpc10nz==7'd123/*US*/))  xpc10nz <= 7'd124/*xpc10nz*/;
                  if ((xpc10nz==7'd124/*US*/))  xpc10nz <= 7'd125/*xpc10nz*/;
                  if ((xpc10nz==7'd125/*US*/))  xpc10nz <= 7'd126/*xpc10nz*/;
                  if ((xpc10nz==7'd126/*US*/))  xpc10nz <= 7'd127/*xpc10nz*/;
                  if ((xpc10nz==7'd127/*US*/))  xpc10nz <= 8'd128/*xpc10nz*/;
                  if ((xpc10nz==8'd128/*US*/))  xpc10nz <= 8'd129/*xpc10nz*/;
                  if ((xpc10nz==8'd129/*US*/))  xpc10nz <= 8'd130/*xpc10nz*/;
                  if ((xpc10nz==8'd130/*US*/))  xpc10nz <= 8'd131/*xpc10nz*/;
                  if ((xpc10nz==8'd131/*US*/))  xpc10nz <= 8'd132/*xpc10nz*/;
                  if ((xpc10nz==8'd132/*US*/))  xpc10nz <= 8'd133/*xpc10nz*/;
                  if ((xpc10nz==8'd133/*US*/))  xpc10nz <= 8'd134/*xpc10nz*/;
                  if ((xpc10nz==8'd134/*US*/))  xpc10nz <= 8'd135/*xpc10nz*/;
                  if ((xpc10nz==8'd135/*US*/))  xpc10nz <= 8'd136/*xpc10nz*/;
                  if ((xpc10nz==8'd136/*US*/))  xpc10nz <= 8'd137/*xpc10nz*/;
                  if ((xpc10nz==8'd137/*US*/))  xpc10nz <= 8'd138/*xpc10nz*/;
                  if ((xpc10nz==8'd138/*US*/))  xpc10nz <= 8'd139/*xpc10nz*/;
                  if ((xpc10nz==8'd139/*US*/))  xpc10nz <= 8'd140/*xpc10nz*/;
                  if ((xpc10nz==8'd140/*US*/))  xpc10nz <= 8'd141/*xpc10nz*/;
                  if ((xpc10nz==8'd141/*US*/))  xpc10nz <= 8'd142/*xpc10nz*/;
                  if ((xpc10nz==8'd142/*US*/))  xpc10nz <= 8'd143/*xpc10nz*/;
                  if ((xpc10nz==8'd143/*US*/))  xpc10nz <= 8'd144/*xpc10nz*/;
                  if ((xpc10nz==8'd144/*US*/))  xpc10nz <= 8'd145/*xpc10nz*/;
                  if ((xpc10nz==8'd145/*US*/))  xpc10nz <= 8'd146/*xpc10nz*/;
                  if ((xpc10nz==8'd146/*US*/))  xpc10nz <= 8'd147/*xpc10nz*/;
                  if ((xpc10nz==8'd147/*US*/))  xpc10nz <= 8'd148/*xpc10nz*/;
                  if ((xpc10nz==8'd148/*US*/))  xpc10nz <= 8'd149/*xpc10nz*/;
                  if ((xpc10nz==8'd149/*US*/))  xpc10nz <= 8'd150/*xpc10nz*/;
                  if ((xpc10nz==8'd150/*US*/))  xpc10nz <= 8'd151/*xpc10nz*/;
                  if ((xpc10nz==8'd151/*US*/))  xpc10nz <= 8'd152/*xpc10nz*/;
                  if ((xpc10nz==8'd152/*US*/))  xpc10nz <= 8'd153/*xpc10nz*/;
                  if ((xpc10nz==8'd153/*US*/))  xpc10nz <= 8'd154/*xpc10nz*/;
                  if ((xpc10nz==8'd154/*US*/))  xpc10nz <= 8'd155/*xpc10nz*/;
                  if ((xpc10nz==8'd155/*US*/))  xpc10nz <= 8'd156/*xpc10nz*/;
                  if ((xpc10nz==8'd156/*US*/))  xpc10nz <= 8'd157/*xpc10nz*/;
                  if ((xpc10nz==8'd157/*US*/))  xpc10nz <= 8'd158/*xpc10nz*/;
                  if ((xpc10nz==8'd158/*US*/))  xpc10nz <= 8'd159/*xpc10nz*/;
                  if ((xpc10nz==8'd159/*US*/))  xpc10nz <= 8'd160/*xpc10nz*/;
                  if ((xpc10nz==8'd160/*US*/))  xpc10nz <= 8'd161/*xpc10nz*/;
                  if ((xpc10nz==8'd161/*US*/))  xpc10nz <= 8'd162/*xpc10nz*/;
                  if ((xpc10nz==8'd162/*US*/))  xpc10nz <= 8'd163/*xpc10nz*/;
                  if ((xpc10nz==8'd163/*US*/))  xpc10nz <= 8'd164/*xpc10nz*/;
                  if ((xpc10nz==8'd164/*US*/))  xpc10nz <= 8'd165/*xpc10nz*/;
                  if ((xpc10nz==8'd165/*US*/))  xpc10nz <= 8'd166/*xpc10nz*/;
                  if ((xpc10nz==8'd166/*US*/))  xpc10nz <= 8'd167/*xpc10nz*/;
                  if ((xpc10nz==8'd167/*US*/))  xpc10nz <= 8'd168/*xpc10nz*/;
                  if ((xpc10nz==8'd168/*US*/))  xpc10nz <= 8'd169/*xpc10nz*/;
                  if ((xpc10nz==8'd169/*US*/))  xpc10nz <= 8'd170/*xpc10nz*/;
                  if ((xpc10nz==8'd172/*US*/))  xpc10nz <= 8'd173/*xpc10nz*/;
                  if ((xpc10nz==8'd173/*US*/))  xpc10nz <= 8'd174/*xpc10nz*/;
                  if ((xpc10nz==8'd174/*US*/))  xpc10nz <= 8'd175/*xpc10nz*/;
                  if ((xpc10nz==8'd175/*US*/))  xpc10nz <= 8'd176/*xpc10nz*/;
                  if ((xpc10nz==8'd176/*US*/))  xpc10nz <= 8'd177/*xpc10nz*/;
                  if ((xpc10nz==8'd177/*US*/))  xpc10nz <= 8'd178/*xpc10nz*/;
                  if ((xpc10nz==8'd178/*US*/))  xpc10nz <= 8'd179/*xpc10nz*/;
                  if ((xpc10nz==8'd179/*US*/))  xpc10nz <= 8'd180/*xpc10nz*/;
                  if ((xpc10nz==8'd180/*US*/))  xpc10nz <= 8'd181/*xpc10nz*/;
                  if ((xpc10nz==8'd181/*US*/))  xpc10nz <= 8'd182/*xpc10nz*/;
                  if ((xpc10nz==8'd182/*US*/))  xpc10nz <= 8'd183/*xpc10nz*/;
                  if ((xpc10nz==8'd183/*US*/))  xpc10nz <= 8'd184/*xpc10nz*/;
                  if ((xpc10nz==8'd184/*US*/))  xpc10nz <= 8'd185/*xpc10nz*/;
                  if ((xpc10nz==8'd185/*US*/))  xpc10nz <= 8'd186/*xpc10nz*/;
                  if ((xpc10nz==8'd186/*US*/))  xpc10nz <= 8'd187/*xpc10nz*/;
                  if ((xpc10nz==8'd187/*US*/))  xpc10nz <= 8'd188/*xpc10nz*/;
                  if ((xpc10nz==8'd188/*US*/))  xpc10nz <= 8'd189/*xpc10nz*/;
                  if ((xpc10nz==8'd189/*US*/))  xpc10nz <= 8'd190/*xpc10nz*/;
                  if ((xpc10nz==8'd190/*US*/))  xpc10nz <= 8'd191/*xpc10nz*/;
                  if ((xpc10nz==8'd191/*US*/))  xpc10nz <= 8'd192/*xpc10nz*/;
                  if ((xpc10nz==8'd192/*US*/))  xpc10nz <= 8'd193/*xpc10nz*/;
                  if ((xpc10nz==8'd193/*US*/))  xpc10nz <= 8'd194/*xpc10nz*/;
                  if ((xpc10nz==8'd194/*US*/))  xpc10nz <= 8'd195/*xpc10nz*/;
                  if ((xpc10nz==8'd195/*US*/))  xpc10nz <= 8'd196/*xpc10nz*/;
                  if ((xpc10nz==8'd196/*US*/))  xpc10nz <= 8'd197/*xpc10nz*/;
                  if ((xpc10nz==8'd197/*US*/))  xpc10nz <= 8'd198/*xpc10nz*/;
                  if ((xpc10nz==8'd198/*US*/))  xpc10nz <= 8'd199/*xpc10nz*/;
                  if ((xpc10nz==8'd199/*US*/))  xpc10nz <= 8'd200/*xpc10nz*/;
                  if ((xpc10nz==8'd200/*US*/))  xpc10nz <= 8'd201/*xpc10nz*/;
                  if ((xpc10nz==8'd201/*US*/))  xpc10nz <= 8'd202/*xpc10nz*/;
                  if ((xpc10nz==8'd202/*US*/))  xpc10nz <= 8'd203/*xpc10nz*/;
                  if ((xpc10nz==8'd203/*US*/))  xpc10nz <= 8'd204/*xpc10nz*/;
                  if ((xpc10nz==8'd204/*US*/))  xpc10nz <= 8'd205/*xpc10nz*/;
                  if ((xpc10nz==8'd205/*US*/))  xpc10nz <= 8'd206/*xpc10nz*/;
                  if ((xpc10nz==8'd206/*US*/))  xpc10nz <= 8'd207/*xpc10nz*/;
                  if ((xpc10nz==8'd207/*US*/))  xpc10nz <= 8'd208/*xpc10nz*/;
                  if ((xpc10nz==8'd208/*US*/))  xpc10nz <= 8'd209/*xpc10nz*/;
                  if ((xpc10nz==8'd209/*US*/))  xpc10nz <= 8'd210/*xpc10nz*/;
                  if ((xpc10nz==8'd210/*US*/))  xpc10nz <= 8'd211/*xpc10nz*/;
                  if ((xpc10nz==8'd211/*US*/))  xpc10nz <= 8'd212/*xpc10nz*/;
                  if ((xpc10nz==8'd212/*US*/))  xpc10nz <= 8'd213/*xpc10nz*/;
                  if ((xpc10nz==8'd213/*US*/))  xpc10nz <= 8'd214/*xpc10nz*/;
                  if ((xpc10nz==8'd214/*US*/))  xpc10nz <= 8'd215/*xpc10nz*/;
                  if ((xpc10nz==8'd215/*US*/))  xpc10nz <= 8'd216/*xpc10nz*/;
                  if ((xpc10nz==8'd216/*US*/))  xpc10nz <= 8'd217/*xpc10nz*/;
                  if ((xpc10nz==8'd217/*US*/))  xpc10nz <= 8'd218/*xpc10nz*/;
                  if ((xpc10nz==8'd218/*US*/))  xpc10nz <= 8'd219/*xpc10nz*/;
                  if ((xpc10nz==8'd219/*US*/))  xpc10nz <= 8'd220/*xpc10nz*/;
                  if ((xpc10nz==8'd220/*US*/))  xpc10nz <= 8'd221/*xpc10nz*/;
                  if ((xpc10nz==8'd221/*US*/))  xpc10nz <= 8'd222/*xpc10nz*/;
                  if ((xpc10nz==8'd222/*US*/))  xpc10nz <= 8'd223/*xpc10nz*/;
                  if ((xpc10nz==8'd223/*US*/))  xpc10nz <= 8'd224/*xpc10nz*/;
                  if ((xpc10nz==8'd224/*US*/))  xpc10nz <= 8'd225/*xpc10nz*/;
                  if ((xpc10nz==8'd225/*US*/))  xpc10nz <= 8'd226/*xpc10nz*/;
                  if ((xpc10nz==8'd226/*US*/))  xpc10nz <= 8'd227/*xpc10nz*/;
                  if ((xpc10nz==8'd227/*US*/))  xpc10nz <= 8'd228/*xpc10nz*/;
                  if ((xpc10nz==8'd228/*US*/))  xpc10nz <= 8'd229/*xpc10nz*/;
                  if ((xpc10nz==8'd229/*US*/))  xpc10nz <= 8'd230/*xpc10nz*/;
                  if ((xpc10nz==8'd230/*US*/))  xpc10nz <= 8'd231/*xpc10nz*/;
                  if ((xpc10nz==8'd231/*US*/))  xpc10nz <= 8'd232/*xpc10nz*/;
                  if ((xpc10nz==8'd232/*US*/))  xpc10nz <= 8'd233/*xpc10nz*/;
                  if ((xpc10nz==8'd233/*US*/))  xpc10nz <= 8'd234/*xpc10nz*/;
                  if ((xpc10nz==8'd234/*US*/))  xpc10nz <= 8'd235/*xpc10nz*/;
                  if ((xpc10nz==8'd236/*US*/))  xpc10nz <= 8'd237/*xpc10nz*/;
                  if ((xpc10nz==8'd239/*US*/))  xpc10nz <= 8'd240/*xpc10nz*/;
                  if ((xpc10nz==9'd256/*US*/))  xpc10nz <= 9'd257/*xpc10nz*/;
                  if ((xpc10nz==9'd260/*US*/))  xpc10nz <= 9'd330/*xpc10nz*/;
                  if ((xpc10nz==9'd261/*US*/))  xpc10nz <= 9'd335/*xpc10nz*/;
                  if ((xpc10nz==9'd262/*US*/))  xpc10nz <= 9'd338/*xpc10nz*/;
                  if ((xpc10nz==9'd263/*US*/))  xpc10nz <= 9'd340/*xpc10nz*/;
                  if ((xpc10nz==9'd264/*US*/))  xpc10nz <= 9'd334/*xpc10nz*/;
                  if ((xpc10nz==9'd265/*US*/))  xpc10nz <= 9'd330/*xpc10nz*/;
                  if ((xpc10nz==9'd266/*US*/))  xpc10nz <= 9'd335/*xpc10nz*/;
                  if ((xpc10nz==9'd267/*US*/))  xpc10nz <= 9'd338/*xpc10nz*/;
                  if ((xpc10nz==9'd268/*US*/))  xpc10nz <= 9'd340/*xpc10nz*/;
                  if ((xpc10nz==9'd269/*US*/))  xpc10nz <= 9'd334/*xpc10nz*/;
                  if ((xpc10nz==9'd270/*US*/))  xpc10nz <= 9'd330/*xpc10nz*/;
                  if ((xpc10nz==9'd271/*US*/))  xpc10nz <= 9'd335/*xpc10nz*/;
                  if ((xpc10nz==9'd272/*US*/))  xpc10nz <= 9'd338/*xpc10nz*/;
                  if ((xpc10nz==9'd273/*US*/))  xpc10nz <= 9'd340/*xpc10nz*/;
                  if ((xpc10nz==9'd274/*US*/))  xpc10nz <= 9'd334/*xpc10nz*/;
                  if ((xpc10nz==9'd275/*US*/))  xpc10nz <= 9'd330/*xpc10nz*/;
                  if ((xpc10nz==9'd276/*US*/))  xpc10nz <= 9'd335/*xpc10nz*/;
                  if ((xpc10nz==9'd277/*US*/))  xpc10nz <= 9'd338/*xpc10nz*/;
                  if ((xpc10nz==9'd278/*US*/))  xpc10nz <= 9'd340/*xpc10nz*/;
                  if ((xpc10nz==9'd279/*US*/))  xpc10nz <= 9'd334/*xpc10nz*/;
                  if ((xpc10nz==9'd280/*US*/))  xpc10nz <= 9'd334/*xpc10nz*/;
                  if ((xpc10nz==9'd281/*US*/))  xpc10nz <= 9'd334/*xpc10nz*/;
                  if ((xpc10nz==9'd282/*US*/))  xpc10nz <= 9'd334/*xpc10nz*/;
                  if ((xpc10nz==9'd283/*US*/))  xpc10nz <= 9'd334/*xpc10nz*/;
                  if ((xpc10nz==9'd285/*US*/))  xpc10nz <= 9'd286/*xpc10nz*/;
                  if ((xpc10nz==9'd287/*US*/))  xpc10nz <= 9'd288/*xpc10nz*/;
                  if ((xpc10nz==9'd290/*US*/))  xpc10nz <= 9'd314/*xpc10nz*/;
                  if ((xpc10nz==9'd291/*US*/))  xpc10nz <= 9'd324/*xpc10nz*/;
                  if ((xpc10nz==9'd292/*US*/))  xpc10nz <= 9'd327/*xpc10nz*/;
                  if ((xpc10nz==9'd293/*US*/))  xpc10nz <= 9'd329/*xpc10nz*/;
                  if ((xpc10nz==9'd294/*US*/))  xpc10nz <= 9'd318/*xpc10nz*/;
                  if ((xpc10nz==9'd295/*US*/))  xpc10nz <= 9'd314/*xpc10nz*/;
                  if ((xpc10nz==9'd296/*US*/))  xpc10nz <= 9'd324/*xpc10nz*/;
                  if ((xpc10nz==9'd297/*US*/))  xpc10nz <= 9'd327/*xpc10nz*/;
                  if ((xpc10nz==9'd298/*US*/))  xpc10nz <= 9'd329/*xpc10nz*/;
                  if ((xpc10nz==9'd299/*US*/))  xpc10nz <= 9'd318/*xpc10nz*/;
                  if ((xpc10nz==9'd300/*US*/))  xpc10nz <= 9'd314/*xpc10nz*/;
                  if ((xpc10nz==9'd301/*US*/))  xpc10nz <= 9'd324/*xpc10nz*/;
                  if ((xpc10nz==9'd302/*US*/))  xpc10nz <= 9'd327/*xpc10nz*/;
                  if ((xpc10nz==9'd303/*US*/))  xpc10nz <= 9'd329/*xpc10nz*/;
                  if ((xpc10nz==9'd304/*US*/))  xpc10nz <= 9'd318/*xpc10nz*/;
                  if ((xpc10nz==9'd305/*US*/))  xpc10nz <= 9'd314/*xpc10nz*/;
                  if ((xpc10nz==9'd306/*US*/))  xpc10nz <= 9'd324/*xpc10nz*/;
                  if ((xpc10nz==9'd307/*US*/))  xpc10nz <= 9'd327/*xpc10nz*/;
                  if ((xpc10nz==9'd308/*US*/))  xpc10nz <= 9'd329/*xpc10nz*/;
                  if ((xpc10nz==9'd309/*US*/))  xpc10nz <= 9'd318/*xpc10nz*/;
                  if ((xpc10nz==9'd310/*US*/))  xpc10nz <= 9'd318/*xpc10nz*/;
                  if ((xpc10nz==9'd311/*US*/))  xpc10nz <= 9'd318/*xpc10nz*/;
                  if ((xpc10nz==9'd312/*US*/))  xpc10nz <= 9'd318/*xpc10nz*/;
                  if ((xpc10nz==9'd313/*US*/))  xpc10nz <= 9'd318/*xpc10nz*/;
                  if ((xpc10nz==9'd315/*US*/))  xpc10nz <= 9'd318/*xpc10nz*/;
                  if ((xpc10nz==9'd316/*US*/))  xpc10nz <= 9'd318/*xpc10nz*/;
                  if ((xpc10nz==9'd317/*US*/))  xpc10nz <= 9'd318/*xpc10nz*/;
                  if ((xpc10nz==9'd325/*US*/))  xpc10nz <= 9'd318/*xpc10nz*/;
                  if ((xpc10nz==9'd326/*US*/))  xpc10nz <= 9'd318/*xpc10nz*/;
                  if ((xpc10nz==9'd328/*US*/))  xpc10nz <= 9'd318/*xpc10nz*/;
                  if ((xpc10nz==9'd331/*US*/))  xpc10nz <= 9'd334/*xpc10nz*/;
                  if ((xpc10nz==9'd332/*US*/))  xpc10nz <= 9'd334/*xpc10nz*/;
                  if ((xpc10nz==9'd333/*US*/))  xpc10nz <= 9'd334/*xpc10nz*/;
                  if ((xpc10nz==9'd336/*US*/))  xpc10nz <= 9'd334/*xpc10nz*/;
                  if ((xpc10nz==9'd337/*US*/))  xpc10nz <= 9'd334/*xpc10nz*/;
                  if ((xpc10nz==9'd339/*US*/))  xpc10nz <= 9'd334/*xpc10nz*/;
                  if ((xpc10nz==9'd343/*US*/))  xpc10nz <= 9'd344/*xpc10nz*/;
                  if ((xpc10nz==9'd344/*US*/))  xpc10nz <= 9'd345/*xpc10nz*/;
                  if ((xpc10nz==9'd345/*US*/))  xpc10nz <= 9'd346/*xpc10nz*/;
                  if ((xpc10nz==9'd346/*US*/))  xpc10nz <= 9'd347/*xpc10nz*/;
                  if ((xpc10nz==9'd347/*US*/))  xpc10nz <= 9'd348/*xpc10nz*/;
                  if ((xpc10nz==9'd348/*US*/))  xpc10nz <= 9'd349/*xpc10nz*/;
                  if ((xpc10nz==9'd349/*US*/))  xpc10nz <= 9'd350/*xpc10nz*/;
                  if ((xpc10nz==9'd350/*US*/))  xpc10nz <= 9'd351/*xpc10nz*/;
                  if ((xpc10nz==9'd351/*US*/))  xpc10nz <= 9'd352/*xpc10nz*/;
                  if ((xpc10nz==9'd352/*US*/))  xpc10nz <= 9'd353/*xpc10nz*/;
                  if ((xpc10nz==9'd353/*US*/))  xpc10nz <= 9'd354/*xpc10nz*/;
                  if ((xpc10nz==9'd354/*US*/))  xpc10nz <= 9'd355/*xpc10nz*/;
                  if ((xpc10nz==9'd355/*US*/))  xpc10nz <= 9'd356/*xpc10nz*/;
                  if ((xpc10nz==9'd356/*US*/))  xpc10nz <= 9'd357/*xpc10nz*/;
                  if ((xpc10nz==9'd357/*US*/))  xpc10nz <= 9'd358/*xpc10nz*/;
                  if ((xpc10nz==9'd358/*US*/))  xpc10nz <= 9'd359/*xpc10nz*/;
                  if ((xpc10nz==9'd359/*US*/))  xpc10nz <= 9'd360/*xpc10nz*/;
                  if ((xpc10nz==9'd360/*US*/))  xpc10nz <= 9'd361/*xpc10nz*/;
                  if ((xpc10nz==9'd361/*US*/))  xpc10nz <= 9'd362/*xpc10nz*/;
                  if ((xpc10nz==9'd362/*US*/))  xpc10nz <= 9'd363/*xpc10nz*/;
                  if ((xpc10nz==9'd363/*US*/))  xpc10nz <= 9'd364/*xpc10nz*/;
                  if ((xpc10nz==9'd364/*US*/))  xpc10nz <= 9'd365/*xpc10nz*/;
                  if ((xpc10nz==9'd365/*US*/))  xpc10nz <= 9'd366/*xpc10nz*/;
                  if ((xpc10nz==9'd366/*US*/))  xpc10nz <= 9'd367/*xpc10nz*/;
                  if ((xpc10nz==9'd367/*US*/))  xpc10nz <= 9'd368/*xpc10nz*/;
                  if ((xpc10nz==9'd368/*US*/))  xpc10nz <= 9'd369/*xpc10nz*/;
                  if ((xpc10nz==9'd369/*US*/))  xpc10nz <= 9'd370/*xpc10nz*/;
                  if ((xpc10nz==9'd370/*US*/))  xpc10nz <= 9'd371/*xpc10nz*/;
                  if ((xpc10nz==9'd371/*US*/))  xpc10nz <= 9'd372/*xpc10nz*/;
                  if ((xpc10nz==9'd372/*US*/))  xpc10nz <= 9'd373/*xpc10nz*/;
                  if ((xpc10nz==9'd373/*US*/))  xpc10nz <= 9'd374/*xpc10nz*/;
                  if ((xpc10nz==9'd374/*US*/))  xpc10nz <= 9'd375/*xpc10nz*/;
                  if ((xpc10nz==9'd375/*US*/))  xpc10nz <= 9'd376/*xpc10nz*/;
                  if ((xpc10nz==9'd376/*US*/))  xpc10nz <= 9'd377/*xpc10nz*/;
                  if ((xpc10nz==9'd377/*US*/))  xpc10nz <= 9'd378/*xpc10nz*/;
                  if ((xpc10nz==9'd378/*US*/))  xpc10nz <= 9'd379/*xpc10nz*/;
                  if ((xpc10nz==9'd379/*US*/))  xpc10nz <= 9'd380/*xpc10nz*/;
                  if ((xpc10nz==9'd380/*US*/))  xpc10nz <= 9'd381/*xpc10nz*/;
                  if ((xpc10nz==9'd381/*US*/))  xpc10nz <= 9'd382/*xpc10nz*/;
                  if ((xpc10nz==9'd382/*US*/))  xpc10nz <= 9'd383/*xpc10nz*/;
                  if ((xpc10nz==9'd383/*US*/))  xpc10nz <= 9'd384/*xpc10nz*/;
                  if ((xpc10nz==9'd384/*US*/))  xpc10nz <= 9'd385/*xpc10nz*/;
                  if ((xpc10nz==9'd385/*US*/))  xpc10nz <= 9'd386/*xpc10nz*/;
                  if ((xpc10nz==9'd386/*US*/))  xpc10nz <= 9'd387/*xpc10nz*/;
                  if ((xpc10nz==9'd387/*US*/))  xpc10nz <= 9'd388/*xpc10nz*/;
                  if ((xpc10nz==9'd388/*US*/))  xpc10nz <= 9'd389/*xpc10nz*/;
                  if ((xpc10nz==9'd389/*US*/))  xpc10nz <= 9'd390/*xpc10nz*/;
                  if ((xpc10nz==9'd390/*US*/))  xpc10nz <= 9'd391/*xpc10nz*/;
                  if ((xpc10nz==9'd391/*US*/))  xpc10nz <= 9'd392/*xpc10nz*/;
                  if ((xpc10nz==9'd392/*US*/))  xpc10nz <= 9'd393/*xpc10nz*/;
                  if ((xpc10nz==9'd393/*US*/))  xpc10nz <= 9'd394/*xpc10nz*/;
                  if ((xpc10nz==9'd394/*US*/))  xpc10nz <= 9'd395/*xpc10nz*/;
                  if ((xpc10nz==9'd395/*US*/))  xpc10nz <= 9'd396/*xpc10nz*/;
                  if ((xpc10nz==9'd396/*US*/))  xpc10nz <= 9'd397/*xpc10nz*/;
                  if ((xpc10nz==9'd397/*US*/))  xpc10nz <= 9'd398/*xpc10nz*/;
                  if ((xpc10nz==9'd398/*US*/))  xpc10nz <= 9'd399/*xpc10nz*/;
                  if ((xpc10nz==9'd399/*US*/))  xpc10nz <= 9'd400/*xpc10nz*/;
                  if ((xpc10nz==9'd400/*US*/))  xpc10nz <= 9'd401/*xpc10nz*/;
                  if ((xpc10nz==9'd401/*US*/))  xpc10nz <= 9'd402/*xpc10nz*/;
                  if ((xpc10nz==9'd402/*US*/))  xpc10nz <= 9'd403/*xpc10nz*/;
                  if ((xpc10nz==9'd403/*US*/))  xpc10nz <= 9'd404/*xpc10nz*/;
                  if ((xpc10nz==9'd404/*US*/))  xpc10nz <= 9'd405/*xpc10nz*/;
                  if ((xpc10nz==9'd405/*US*/))  xpc10nz <= 9'd406/*xpc10nz*/;
                  if ((xpc10nz==9'd408/*US*/))  xpc10nz <= 9'd409/*xpc10nz*/;
                  if ((xpc10nz==9'd409/*US*/))  xpc10nz <= 9'd410/*xpc10nz*/;
                  if ((xpc10nz==9'd410/*US*/))  xpc10nz <= 9'd411/*xpc10nz*/;
                  if ((xpc10nz==9'd411/*US*/))  xpc10nz <= 9'd412/*xpc10nz*/;
                  if ((xpc10nz==9'd412/*US*/))  xpc10nz <= 9'd413/*xpc10nz*/;
                  if ((xpc10nz==9'd413/*US*/))  xpc10nz <= 9'd414/*xpc10nz*/;
                  if ((xpc10nz==9'd414/*US*/))  xpc10nz <= 9'd415/*xpc10nz*/;
                  if ((xpc10nz==9'd415/*US*/))  xpc10nz <= 9'd416/*xpc10nz*/;
                  if ((xpc10nz==9'd416/*US*/))  xpc10nz <= 9'd417/*xpc10nz*/;
                  if ((xpc10nz==9'd417/*US*/))  xpc10nz <= 9'd418/*xpc10nz*/;
                  if ((xpc10nz==9'd418/*US*/))  xpc10nz <= 9'd419/*xpc10nz*/;
                  if ((xpc10nz==9'd419/*US*/))  xpc10nz <= 9'd420/*xpc10nz*/;
                  if ((xpc10nz==9'd420/*US*/))  xpc10nz <= 9'd421/*xpc10nz*/;
                  if ((xpc10nz==9'd421/*US*/))  xpc10nz <= 9'd422/*xpc10nz*/;
                  if ((xpc10nz==9'd422/*US*/))  xpc10nz <= 9'd423/*xpc10nz*/;
                  if ((xpc10nz==9'd423/*US*/))  xpc10nz <= 9'd424/*xpc10nz*/;
                  if ((xpc10nz==9'd424/*US*/))  xpc10nz <= 9'd425/*xpc10nz*/;
                  if ((xpc10nz==9'd425/*US*/))  xpc10nz <= 9'd426/*xpc10nz*/;
                  if ((xpc10nz==9'd426/*US*/))  xpc10nz <= 9'd427/*xpc10nz*/;
                  if ((xpc10nz==9'd427/*US*/))  xpc10nz <= 9'd428/*xpc10nz*/;
                  if ((xpc10nz==9'd428/*US*/))  xpc10nz <= 9'd429/*xpc10nz*/;
                  if ((xpc10nz==9'd429/*US*/))  xpc10nz <= 9'd430/*xpc10nz*/;
                  if ((xpc10nz==9'd430/*US*/))  xpc10nz <= 9'd431/*xpc10nz*/;
                  if ((xpc10nz==9'd431/*US*/))  xpc10nz <= 9'd432/*xpc10nz*/;
                  if ((xpc10nz==9'd432/*US*/))  xpc10nz <= 9'd433/*xpc10nz*/;
                  if ((xpc10nz==9'd433/*US*/))  xpc10nz <= 9'd434/*xpc10nz*/;
                  if ((xpc10nz==9'd434/*US*/))  xpc10nz <= 9'd435/*xpc10nz*/;
                  if ((xpc10nz==9'd435/*US*/))  xpc10nz <= 9'd436/*xpc10nz*/;
                  if ((xpc10nz==9'd436/*US*/))  xpc10nz <= 9'd437/*xpc10nz*/;
                  if ((xpc10nz==9'd437/*US*/))  xpc10nz <= 9'd438/*xpc10nz*/;
                  if ((xpc10nz==9'd438/*US*/))  xpc10nz <= 9'd439/*xpc10nz*/;
                  if ((xpc10nz==9'd439/*US*/))  xpc10nz <= 9'd440/*xpc10nz*/;
                  if ((xpc10nz==9'd440/*US*/))  xpc10nz <= 9'd441/*xpc10nz*/;
                  if ((xpc10nz==9'd441/*US*/))  xpc10nz <= 9'd442/*xpc10nz*/;
                  if ((xpc10nz==9'd442/*US*/))  xpc10nz <= 9'd443/*xpc10nz*/;
                  if ((xpc10nz==9'd443/*US*/))  xpc10nz <= 9'd444/*xpc10nz*/;
                  if ((xpc10nz==9'd444/*US*/))  xpc10nz <= 9'd445/*xpc10nz*/;
                  if ((xpc10nz==9'd445/*US*/))  xpc10nz <= 9'd446/*xpc10nz*/;
                  if ((xpc10nz==9'd446/*US*/))  xpc10nz <= 9'd447/*xpc10nz*/;
                  if ((xpc10nz==9'd447/*US*/))  xpc10nz <= 9'd448/*xpc10nz*/;
                  if ((xpc10nz==9'd448/*US*/))  xpc10nz <= 9'd449/*xpc10nz*/;
                  if ((xpc10nz==9'd449/*US*/))  xpc10nz <= 9'd450/*xpc10nz*/;
                  if ((xpc10nz==9'd450/*US*/))  xpc10nz <= 9'd451/*xpc10nz*/;
                  if ((xpc10nz==9'd451/*US*/))  xpc10nz <= 9'd452/*xpc10nz*/;
                  if ((xpc10nz==9'd452/*US*/))  xpc10nz <= 9'd453/*xpc10nz*/;
                  if ((xpc10nz==9'd453/*US*/))  xpc10nz <= 9'd454/*xpc10nz*/;
                  if ((xpc10nz==9'd454/*US*/))  xpc10nz <= 9'd455/*xpc10nz*/;
                  if ((xpc10nz==9'd455/*US*/))  xpc10nz <= 9'd456/*xpc10nz*/;
                  if ((xpc10nz==9'd456/*US*/))  xpc10nz <= 9'd457/*xpc10nz*/;
                  if ((xpc10nz==9'd457/*US*/))  xpc10nz <= 9'd458/*xpc10nz*/;
                  if ((xpc10nz==9'd458/*US*/))  xpc10nz <= 9'd459/*xpc10nz*/;
                  if ((xpc10nz==9'd459/*US*/))  xpc10nz <= 9'd460/*xpc10nz*/;
                  if ((xpc10nz==9'd460/*US*/))  xpc10nz <= 9'd461/*xpc10nz*/;
                  if ((xpc10nz==9'd461/*US*/))  xpc10nz <= 9'd462/*xpc10nz*/;
                  if ((xpc10nz==9'd462/*US*/))  xpc10nz <= 9'd463/*xpc10nz*/;
                  if ((xpc10nz==9'd463/*US*/))  xpc10nz <= 9'd464/*xpc10nz*/;
                  if ((xpc10nz==9'd464/*US*/))  xpc10nz <= 9'd465/*xpc10nz*/;
                  if ((xpc10nz==9'd465/*US*/))  xpc10nz <= 9'd466/*xpc10nz*/;
                  if ((xpc10nz==9'd466/*US*/))  xpc10nz <= 9'd467/*xpc10nz*/;
                  if ((xpc10nz==9'd467/*US*/))  xpc10nz <= 9'd468/*xpc10nz*/;
                  if ((xpc10nz==9'd468/*US*/))  xpc10nz <= 9'd469/*xpc10nz*/;
                  if ((xpc10nz==9'd469/*US*/))  xpc10nz <= 9'd470/*xpc10nz*/;
                  if ((xpc10nz==9'd470/*US*/))  xpc10nz <= 9'd471/*xpc10nz*/;
                  if ((xpc10nz==9'd472/*US*/))  xpc10nz <= 9'd473/*xpc10nz*/;
                  if ((xpc10nz==9'd474/*US*/))  xpc10nz <= 9'd502/*xpc10nz*/;
                  if ((xpc10nz==9'd475/*US*/))  xpc10nz <= 9'd330/*xpc10nz*/;
                  if ((xpc10nz==9'd476/*US*/))  xpc10nz <= 9'd335/*xpc10nz*/;
                  if ((xpc10nz==9'd477/*US*/))  xpc10nz <= 9'd338/*xpc10nz*/;
                  if ((xpc10nz==9'd478/*US*/))  xpc10nz <= 9'd340/*xpc10nz*/;
                  if ((xpc10nz==9'd479/*US*/))  xpc10nz <= 9'd334/*xpc10nz*/;
                  if ((xpc10nz==9'd480/*US*/))  xpc10nz <= 9'd502/*xpc10nz*/;
                  if ((xpc10nz==9'd481/*US*/))  xpc10nz <= 9'd330/*xpc10nz*/;
                  if ((xpc10nz==9'd482/*US*/))  xpc10nz <= 9'd335/*xpc10nz*/;
                  if ((xpc10nz==9'd483/*US*/))  xpc10nz <= 9'd338/*xpc10nz*/;
                  if ((xpc10nz==9'd484/*US*/))  xpc10nz <= 9'd340/*xpc10nz*/;
                  if ((xpc10nz==9'd485/*US*/))  xpc10nz <= 9'd334/*xpc10nz*/;
                  if ((xpc10nz==9'd486/*US*/))  xpc10nz <= 9'd502/*xpc10nz*/;
                  if ((xpc10nz==9'd487/*US*/))  xpc10nz <= 9'd330/*xpc10nz*/;
                  if ((xpc10nz==9'd488/*US*/))  xpc10nz <= 9'd335/*xpc10nz*/;
                  if ((xpc10nz==9'd489/*US*/))  xpc10nz <= 9'd338/*xpc10nz*/;
                  if ((xpc10nz==9'd490/*US*/))  xpc10nz <= 9'd340/*xpc10nz*/;
                  if ((xpc10nz==9'd491/*US*/))  xpc10nz <= 9'd334/*xpc10nz*/;
                  if ((xpc10nz==9'd492/*US*/))  xpc10nz <= 9'd502/*xpc10nz*/;
                  if ((xpc10nz==9'd493/*US*/))  xpc10nz <= 9'd330/*xpc10nz*/;
                  if ((xpc10nz==9'd494/*US*/))  xpc10nz <= 9'd335/*xpc10nz*/;
                  if ((xpc10nz==9'd495/*US*/))  xpc10nz <= 9'd338/*xpc10nz*/;
                  if ((xpc10nz==9'd496/*US*/))  xpc10nz <= 9'd340/*xpc10nz*/;
                  if ((xpc10nz==9'd497/*US*/))  xpc10nz <= 9'd334/*xpc10nz*/;
                  if ((xpc10nz==9'd498/*US*/))  xpc10nz <= 9'd334/*xpc10nz*/;
                  if ((xpc10nz==9'd499/*US*/))  xpc10nz <= 9'd334/*xpc10nz*/;
                  if ((xpc10nz==9'd500/*US*/))  xpc10nz <= 9'd334/*xpc10nz*/;
                  if ((xpc10nz==9'd501/*US*/))  xpc10nz <= 9'd334/*xpc10nz*/;
                  if ((xpc10nz==9'd504/*US*/))  xpc10nz <= 9'd330/*xpc10nz*/;
                  if ((xpc10nz==9'd505/*US*/))  xpc10nz <= 9'd335/*xpc10nz*/;
                  if ((xpc10nz==9'd506/*US*/))  xpc10nz <= 9'd338/*xpc10nz*/;
                  if ((xpc10nz==9'd507/*US*/))  xpc10nz <= 9'd340/*xpc10nz*/;
                  if ((xpc10nz==9'd508/*US*/))  xpc10nz <= 9'd334/*xpc10nz*/;
                  if ((xpc10nz==9'd509/*US*/))  xpc10nz <= 9'd330/*xpc10nz*/;
                  if ((xpc10nz==9'd510/*US*/))  xpc10nz <= 9'd335/*xpc10nz*/;
                  if ((xpc10nz==9'd511/*US*/))  xpc10nz <= 9'd338/*xpc10nz*/;
                  if ((xpc10nz==10'd512/*US*/))  xpc10nz <= 9'd340/*xpc10nz*/;
                  if ((xpc10nz==10'd513/*US*/))  xpc10nz <= 9'd334/*xpc10nz*/;
                  if ((xpc10nz==10'd514/*US*/))  xpc10nz <= 9'd330/*xpc10nz*/;
                  if ((xpc10nz==10'd515/*US*/))  xpc10nz <= 9'd335/*xpc10nz*/;
                  if ((xpc10nz==10'd516/*US*/))  xpc10nz <= 9'd338/*xpc10nz*/;
                  if ((xpc10nz==10'd517/*US*/))  xpc10nz <= 9'd340/*xpc10nz*/;
                  if ((xpc10nz==10'd518/*US*/))  xpc10nz <= 9'd334/*xpc10nz*/;
                  if ((xpc10nz==10'd519/*US*/))  xpc10nz <= 9'd330/*xpc10nz*/;
                  if ((xpc10nz==10'd520/*US*/))  xpc10nz <= 9'd335/*xpc10nz*/;
                  if ((xpc10nz==10'd521/*US*/))  xpc10nz <= 9'd338/*xpc10nz*/;
                  if ((xpc10nz==10'd522/*US*/))  xpc10nz <= 9'd340/*xpc10nz*/;
                  if ((xpc10nz==10'd523/*US*/))  xpc10nz <= 9'd334/*xpc10nz*/;
                  if ((xpc10nz==10'd524/*US*/))  xpc10nz <= 9'd334/*xpc10nz*/;
                  if ((xpc10nz==10'd525/*US*/))  xpc10nz <= 9'd334/*xpc10nz*/;
                  if ((xpc10nz==10'd526/*US*/))  xpc10nz <= 9'd334/*xpc10nz*/;
                  if ((xpc10nz==10'd527/*US*/))  xpc10nz <= 9'd334/*xpc10nz*/;
                  if ((xpc10nz==10'd529/*US*/))  xpc10nz <= 10'd532/*xpc10nz*/;
                  if ((xpc10nz==10'd530/*US*/))  xpc10nz <= 10'd532/*xpc10nz*/;
                  if ((xpc10nz==10'd531/*US*/))  xpc10nz <= 10'd532/*xpc10nz*/;
                  if ((xpc10nz==10'd533/*US*/))  xpc10nz <= 10'd532/*xpc10nz*/;
                  if ((xpc10nz==10'd535/*US*/))  xpc10nz <= 10'd532/*xpc10nz*/;
                  if ((xpc10nz==10'd536/*US*/))  xpc10nz <= 10'd532/*xpc10nz*/;
                  if ((xpc10nz==10'd538/*US*/))  xpc10nz <= 10'd532/*xpc10nz*/;
                  if ((xpc10nz==10'd541/*US*/))  xpc10nz <= 7'd64/*xpc10nz*/;
                  if ((xpc10nz==10'd542/*US*/))  xpc10nz <= 7'd64/*xpc10nz*/;
                  if ((xpc10nz==10'd543/*US*/))  xpc10nz <= 7'd64/*xpc10nz*/;
                  if ((xpc10nz==10'd545/*US*/))  xpc10nz <= 7'd64/*xpc10nz*/;
                  if ((xpc10nz==10'd546/*US*/))  xpc10nz <= 7'd64/*xpc10nz*/;
                  if ((xpc10nz==10'd548/*US*/))  xpc10nz <= 7'd64/*xpc10nz*/;
                  if ((xpc10nz==10'd551/*US*/))  xpc10nz <= 6'd59/*xpc10nz*/;
                  if ((xpc10nz==10'd552/*US*/))  xpc10nz <= 6'd59/*xpc10nz*/;
                  if ((xpc10nz==10'd553/*US*/))  xpc10nz <= 6'd59/*xpc10nz*/;
                  if ((xpc10nz==10'd554/*US*/))  xpc10nz <= 10'd540/*xpc10nz*/;
                  if ((xpc10nz==10'd555/*US*/))  xpc10nz <= 10'd544/*xpc10nz*/;
                  if ((xpc10nz==10'd556/*US*/))  xpc10nz <= 10'd547/*xpc10nz*/;
                  if ((xpc10nz==10'd557/*US*/))  xpc10nz <= 10'd549/*xpc10nz*/;
                  if ((xpc10nz==10'd559/*US*/))  xpc10nz <= 6'd59/*xpc10nz*/;
                  if ((xpc10nz==10'd560/*US*/))  xpc10nz <= 6'd59/*xpc10nz*/;
                  if ((xpc10nz==10'd561/*US*/))  xpc10nz <= 10'd540/*xpc10nz*/;
                  if ((xpc10nz==10'd562/*US*/))  xpc10nz <= 10'd544/*xpc10nz*/;
                  if ((xpc10nz==10'd563/*US*/))  xpc10nz <= 10'd547/*xpc10nz*/;
                  if ((xpc10nz==10'd564/*US*/))  xpc10nz <= 10'd549/*xpc10nz*/;
                  if ((xpc10nz==10'd566/*US*/))  xpc10nz <= 6'd59/*xpc10nz*/;
                  if ((xpc10nz==10'd567/*US*/))  xpc10nz <= 10'd540/*xpc10nz*/;
                  if ((xpc10nz==10'd568/*US*/))  xpc10nz <= 10'd544/*xpc10nz*/;
                  if ((xpc10nz==10'd569/*US*/))  xpc10nz <= 10'd547/*xpc10nz*/;
                  if ((xpc10nz==10'd570/*US*/))  xpc10nz <= 10'd549/*xpc10nz*/;
                  if ((xpc10nz==10'd572/*US*/))  xpc10nz <= 10'd540/*xpc10nz*/;
                  if ((xpc10nz==10'd573/*US*/))  xpc10nz <= 10'd544/*xpc10nz*/;
                  if ((xpc10nz==10'd574/*US*/))  xpc10nz <= 10'd547/*xpc10nz*/;
                  if ((xpc10nz==10'd575/*US*/))  xpc10nz <= 10'd549/*xpc10nz*/;
                  if ((xpc10nz==10'd577/*US*/))  xpc10nz <= 6'd50/*xpc10nz*/;
                  if ((xpc10nz==10'd578/*US*/))  xpc10nz <= 6'd50/*xpc10nz*/;
                  if ((xpc10nz==10'd579/*US*/))  xpc10nz <= 6'd50/*xpc10nz*/;
                  if ((xpc10nz==10'd580/*US*/))  xpc10nz <= 10'd550/*xpc10nz*/;
                  if ((xpc10nz==10'd581/*US*/))  xpc10nz <= 10'd558/*xpc10nz*/;
                  if ((xpc10nz==10'd582/*US*/))  xpc10nz <= 10'd565/*xpc10nz*/;
                  if ((xpc10nz==10'd583/*US*/))  xpc10nz <= 10'd571/*xpc10nz*/;
                  if ((xpc10nz==10'd584/*US*/))  xpc10nz <= 10'd540/*xpc10nz*/;
                  if ((xpc10nz==10'd585/*US*/))  xpc10nz <= 10'd544/*xpc10nz*/;
                  if ((xpc10nz==10'd586/*US*/))  xpc10nz <= 10'd547/*xpc10nz*/;
                  if ((xpc10nz==10'd587/*US*/))  xpc10nz <= 10'd549/*xpc10nz*/;
                  if ((xpc10nz==10'd589/*US*/))  xpc10nz <= 6'd50/*xpc10nz*/;
                  if ((xpc10nz==10'd590/*US*/))  xpc10nz <= 6'd50/*xpc10nz*/;
                  if ((xpc10nz==10'd591/*US*/))  xpc10nz <= 10'd550/*xpc10nz*/;
                  if ((xpc10nz==10'd592/*US*/))  xpc10nz <= 10'd558/*xpc10nz*/;
                  if ((xpc10nz==10'd593/*US*/))  xpc10nz <= 10'd565/*xpc10nz*/;
                  if ((xpc10nz==10'd594/*US*/))  xpc10nz <= 10'd571/*xpc10nz*/;
                  if ((xpc10nz==10'd595/*US*/))  xpc10nz <= 10'd540/*xpc10nz*/;
                  if ((xpc10nz==10'd596/*US*/))  xpc10nz <= 10'd544/*xpc10nz*/;
                  if ((xpc10nz==10'd597/*US*/))  xpc10nz <= 10'd547/*xpc10nz*/;
                  if ((xpc10nz==10'd598/*US*/))  xpc10nz <= 10'd549/*xpc10nz*/;
                  if ((xpc10nz==10'd600/*US*/))  xpc10nz <= 6'd50/*xpc10nz*/;
                  if ((xpc10nz==10'd601/*US*/))  xpc10nz <= 10'd550/*xpc10nz*/;
                  if ((xpc10nz==10'd602/*US*/))  xpc10nz <= 10'd558/*xpc10nz*/;
                  if ((xpc10nz==10'd603/*US*/))  xpc10nz <= 10'd565/*xpc10nz*/;
                  if ((xpc10nz==10'd604/*US*/))  xpc10nz <= 10'd571/*xpc10nz*/;
                  if ((xpc10nz==10'd605/*US*/))  xpc10nz <= 10'd540/*xpc10nz*/;
                  if ((xpc10nz==10'd606/*US*/))  xpc10nz <= 10'd544/*xpc10nz*/;
                  if ((xpc10nz==10'd607/*US*/))  xpc10nz <= 10'd547/*xpc10nz*/;
                  if ((xpc10nz==10'd608/*US*/))  xpc10nz <= 10'd549/*xpc10nz*/;
                  if ((xpc10nz==10'd610/*US*/))  xpc10nz <= 10'd550/*xpc10nz*/;
                  if ((xpc10nz==10'd611/*US*/))  xpc10nz <= 10'd558/*xpc10nz*/;
                  if ((xpc10nz==10'd612/*US*/))  xpc10nz <= 10'd565/*xpc10nz*/;
                  if ((xpc10nz==10'd613/*US*/))  xpc10nz <= 10'd571/*xpc10nz*/;
                  if ((xpc10nz==10'd614/*US*/))  xpc10nz <= 10'd540/*xpc10nz*/;
                  if ((xpc10nz==10'd615/*US*/))  xpc10nz <= 10'd544/*xpc10nz*/;
                  if ((xpc10nz==10'd616/*US*/))  xpc10nz <= 10'd547/*xpc10nz*/;
                  if ((xpc10nz==10'd617/*US*/))  xpc10nz <= 10'd549/*xpc10nz*/;
                   end 
              //End structure HPR cuckoo_hash_demo.exe


       end 
      

  CV_SP_SSRAM_FL1 #(6'd32, 4'd13, 14'd8192, 6'd32) A_SINT_CC_MAPR10NoCE3_ARA0(clk, reset, A_SINT_CC_MAPR10NoCE3_ARA0_RDD0, A_SINT_CC_MAPR10NoCE3_ARA0_AD0
, A_SINT_CC_MAPR10NoCE3_ARA0_WEN0, A_SINT_CC_MAPR10NoCE3_ARA0_REN0, A_SINT_CC_MAPR10NoCE3_ARA0_WRD0);

  CV_SP_SSRAM_FL1 #(6'd32, 4'd13, 14'd8192, 6'd32) A_SINT_CC_MAPR10NoCE2_ARA0(clk, reset, A_SINT_CC_MAPR10NoCE2_ARA0_RDD0, A_SINT_CC_MAPR10NoCE2_ARA0_AD0
, A_SINT_CC_MAPR10NoCE2_ARA0_WEN0, A_SINT_CC_MAPR10NoCE2_ARA0_REN0, A_SINT_CC_MAPR10NoCE2_ARA0_WRD0);

  CV_SP_SSRAM_FL1 #(6'd32, 4'd13, 14'd8192, 6'd32) A_SINT_CC_MAPR10NoCE1_ARA0(clk, reset, A_SINT_CC_MAPR10NoCE1_ARA0_RDD0, A_SINT_CC_MAPR10NoCE1_ARA0_AD0
, A_SINT_CC_MAPR10NoCE1_ARA0_WEN0, A_SINT_CC_MAPR10NoCE1_ARA0_REN0, A_SINT_CC_MAPR10NoCE1_ARA0_WRD0);

  CV_SP_SSRAM_FL1 #(6'd32, 4'd13, 14'd8192, 6'd32) A_SINT_CC_MAPR10NoCE0_ARA0(clk, reset, A_SINT_CC_MAPR10NoCE0_ARA0_RDD0, A_SINT_CC_MAPR10NoCE0_ARA0_AD0
, A_SINT_CC_MAPR10NoCE0_ARA0_WEN0, A_SINT_CC_MAPR10NoCE0_ARA0_REN0, A_SINT_CC_MAPR10NoCE0_ARA0_WRD0);

  CV_INT_VL_MODULUS_S isMODULUS10(clk, reset, isMODULUS10_rdy, isMODULUS10_req, isMODULUS10_RR, isMODULUS10_NN, isMODULUS10_DD, isMODULUS10_err
);

  CV_SP_SSRAM_FL1 #(6'd32, 4'd13, 14'd8192, 6'd32) A_SINT_CC_MAPR12NoCE3_ARB0(clk, reset, A_SINT_CC_MAPR12NoCE3_ARB0_RDD0, A_SINT_CC_MAPR12NoCE3_ARB0_AD0
, A_SINT_CC_MAPR12NoCE3_ARB0_WEN0, A_SINT_CC_MAPR12NoCE3_ARB0_REN0, A_SINT_CC_MAPR12NoCE3_ARB0_WRD0);

  CV_SP_SSRAM_FL1 #(6'd32, 4'd13, 14'd8192, 6'd32) A_SINT_CC_MAPR12NoCE2_ARB0(clk, reset, A_SINT_CC_MAPR12NoCE2_ARB0_RDD0, A_SINT_CC_MAPR12NoCE2_ARB0_AD0
, A_SINT_CC_MAPR12NoCE2_ARB0_WEN0, A_SINT_CC_MAPR12NoCE2_ARB0_REN0, A_SINT_CC_MAPR12NoCE2_ARB0_WRD0);

  CV_SP_SSRAM_FL1 #(6'd32, 4'd13, 14'd8192, 6'd32) A_SINT_CC_MAPR12NoCE1_ARB0(clk, reset, A_SINT_CC_MAPR12NoCE1_ARB0_RDD0, A_SINT_CC_MAPR12NoCE1_ARB0_AD0
, A_SINT_CC_MAPR12NoCE1_ARB0_WEN0, A_SINT_CC_MAPR12NoCE1_ARB0_REN0, A_SINT_CC_MAPR12NoCE1_ARB0_WRD0);

  CV_SP_SSRAM_FL1 #(6'd32, 4'd13, 14'd8192, 6'd32) A_SINT_CC_MAPR12NoCE0_ARB0(clk, reset, A_SINT_CC_MAPR12NoCE0_ARB0_RDD0, A_SINT_CC_MAPR12NoCE0_ARB0_AD0
, A_SINT_CC_MAPR12NoCE0_ARB0_WEN0, A_SINT_CC_MAPR12NoCE0_ARB0_REN0, A_SINT_CC_MAPR12NoCE0_ARB0_WRD0);

  CV_SP_SSRAM_FL1 #(7'd64, 4'd15, 16'd32768, 7'd64) A_64_US_CC_SCALbx26_ARA0(clk, reset, A_64_US_CC_SCALbx26_ARA0_RDD0, A_64_US_CC_SCALbx26_ARA0_AD0
, A_64_US_CC_SCALbx26_ARA0_WEN0, A_64_US_CC_SCALbx26_ARA0_REN0, A_64_US_CC_SCALbx26_ARA0_WRD0);

always @(*) xpc10_clear = (xpc10nz==0/*US*/) || (xpc10nz==1'd1/*US*/) || (xpc10nz==2'd2/*US*/) || (xpc10nz==2'd3/*US*/) || (xpc10nz==3'd4/*US*/) || (xpc10nz==3'd5
/*US*/) || (xpc10nz==3'd6/*US*/) || (xpc10nz==3'd7/*US*/) || (xpc10nz==4'd8/*US*/) || (xpc10nz==4'd9/*US*/) || (xpc10nz==4'd10/*US*/) || 
(xpc10nz==4'd11/*US*/) || (xpc10nz==4'd12/*US*/) || (xpc10nz==4'd13/*US*/) || (xpc10nz==4'd14/*US*/) || (xpc10nz==4'd15/*US*/) || (xpc10nz
==5'd16/*US*/) || (xpc10nz==5'd17/*US*/) || (xpc10nz==5'd18/*US*/) || (xpc10nz==5'd19/*US*/) || (xpc10nz==5'd20/*US*/) || (xpc10nz==6'd37
/*US*/) || (xpc10nz==6'd50/*US*/) || (xpc10nz==6'd59/*US*/) || (xpc10nz==7'd64/*US*/) || (xpc10nz==7'd65/*US*/) || (xpc10nz==7'd82/*US*/) || 
(xpc10nz==7'd83/*US*/) || (xpc10nz==7'd84/*US*/) || (xpc10nz==7'd85/*US*/) || (xpc10nz==7'd86/*US*/) || (xpc10nz==7'd87/*US*/) || (xpc10nz
==7'd88/*US*/) || (xpc10nz==7'd89/*US*/) || (xpc10nz==7'd90/*US*/) || (xpc10nz==7'd91/*US*/) || (xpc10nz==7'd92/*US*/) || (xpc10nz==7'd93
/*US*/) || (xpc10nz==7'd94/*US*/) || (xpc10nz==7'd95/*US*/) || (xpc10nz==7'd96/*US*/) || (xpc10nz==7'd97/*US*/) || (xpc10nz==7'd98/*US*/) || 
(xpc10nz==7'd99/*US*/) || (xpc10nz==7'd100/*US*/) || (xpc10nz==7'd101/*US*/) || (xpc10nz==7'd102/*US*/) || (xpc10nz==7'd103/*US*/) || 
(xpc10nz==7'd104/*US*/) || (xpc10nz==7'd105/*US*/) || (xpc10nz==7'd106/*US*/) || (xpc10nz==8'd171/*US*/) || (xpc10nz==8'd236/*US*/) || 
(xpc10nz==8'd238/*US*/) || (xpc10nz==8'd239/*US*/) || (xpc10nz==8'd241/*US*/) || (xpc10nz==8'd242/*US*/) || (xpc10nz==8'd244/*US*/) || 
(xpc10nz==8'd245/*US*/) || (xpc10nz==8'd246/*US*/) || (xpc10nz==8'd247/*US*/) || (xpc10nz==8'd248/*US*/) || (xpc10nz==8'd249/*US*/) || 
(xpc10nz==8'd250/*US*/) || (xpc10nz==8'd251/*US*/) || (xpc10nz==8'd252/*US*/) || (xpc10nz==8'd253/*US*/) || (xpc10nz==8'd254/*US*/) || 
(xpc10nz==8'd255/*US*/) || (xpc10nz==9'd257/*US*/) || (xpc10nz==9'd258/*US*/) || (xpc10nz==9'd259/*US*/) || (xpc10nz==9'd284/*US*/) || 
(xpc10nz==9'd285/*US*/) || (xpc10nz==9'd287/*US*/) || (xpc10nz==9'd289/*US*/) || (xpc10nz==9'd314/*US*/) || (xpc10nz==9'd318/*US*/) || 
(xpc10nz==9'd319/*US*/) || (xpc10nz==9'd320/*US*/) || (xpc10nz==9'd321/*US*/) || (xpc10nz==9'd322/*US*/) || (xpc10nz==9'd323/*US*/) || 
(xpc10nz==9'd324/*US*/) || (xpc10nz==9'd327/*US*/) || (xpc10nz==9'd329/*US*/) || (xpc10nz==9'd330/*US*/) || (xpc10nz==9'd334/*US*/) || 
(xpc10nz==9'd335/*US*/) || (xpc10nz==9'd338/*US*/) || (xpc10nz==9'd340/*US*/) || (xpc10nz==9'd341/*US*/) || (xpc10nz==9'd342/*US*/) || 
(xpc10nz==9'd407/*US*/) || (xpc10nz==9'd472/*US*/) || (xpc10nz==9'd502/*US*/) || (xpc10nz==9'd503/*US*/) || (xpc10nz==10'd528/*US*/) || 
(xpc10nz==10'd532/*US*/) || (xpc10nz==10'd534/*US*/) || (xpc10nz==10'd537/*US*/) || (xpc10nz==10'd539/*US*/) || (xpc10nz==10'd540/*US*/) || 
(xpc10nz==10'd544/*US*/) || (xpc10nz==10'd547/*US*/) || (xpc10nz==10'd549/*US*/) || (xpc10nz==10'd550/*US*/) || (xpc10nz==10'd558/*US*/) || 
(xpc10nz==10'd565/*US*/) || (xpc10nz==10'd571/*US*/) || (xpc10nz==10'd576/*US*/) || (xpc10nz==10'd588/*US*/) || (xpc10nz==10'd609/*US*/) || 
(xpc10nz==10'd599/*US*/);

always @(*) xpc10_stall = ((xpc10nz==8'd170/*US*/) || (xpc10nz==8'd235/*US*/) || (xpc10nz==9'd406/*US*/) || (xpc10nz==9'd471/*US*/)) && !isMODULUS10_rdy && !isMODULUS10RRh10vld
;

// 1 vectors of width 10
// 28 vectors of width 32
// 97 vectors of width 1
// 10 vectors of width 64
// 1 vectors of width 15
// 8 vectors of width 13
// 8 array locations of width 32
// 928 bits in scalar variables
// Total state bits in module = 2946 bits.
// 354 continuously assigned (wire/non-state) bits 
//   cell CV_SP_SSRAM_FL1 count=9
//   cell CV_INT_VL_MODULUS_S count=1
// Total number of leaf cells = 10
endmodule

//  
// LCP delay estimations included: turn off with -vnl-lcp-delay-estimate=disable
//HPR L/S (orangepath) auxiliary reports.
//KiwiC compilation report
//Kiwi Scientific Acceleration (KiwiC .net/CIL/C# to Verilog/SystemC compiler): Version alpha 2.15f : 19th-June-2016
//22/06/2016 08:19:19
//Cmd line args:  /home/djg11/d320/hprls/kiwipro/kiwic/distro/lib/kiwic.exe -give-backtrace -vnl=cuckoo_hash_demo.v cuckoo_hash_demo.exe -vnl-resets=synchronous -kiwic-cil-dump=combined -kiwic-kcode-dump=enable -res2-loadstore-port-count=0 -vnl-roundtrip=disable -bevelab-default-pause-mode=soft -bevelab-soft-pause-threshold=10 -vnl-rootmodname=DUT


//----------------------------------------------------------

//Report from KiwiC-fe.rpt:::
//KiwiC: front end input processing of class or method called KiwiSystem/Kiwi
//
//root_walk start thread at a static method (used as an entry point). Method name=.cctor uid=cctor10
//
//KiwiC start_thread (or entry point) id=cctor10
//
//Root method elaborated: specificf=S_kickoff_collate leftover=1+0
//
//KiwiC: front end input processing of class or method called System/BitConverter
//
//root_walk start thread at a static method (used as an entry point). Method name=.cctor uid=cctor12
//
//KiwiC start_thread (or entry point) id=cctor12
//
//Root method elaborated: specificf=S_kickoff_collate leftover=1+1
//
//KiwiC: front end input processing of class or method called Testbench
//
//root_walk start thread at a static method (used as an entry point). Method name=.cctor uid=cctor14
//
//KiwiC start_thread (or entry point) id=cctor14
//
//Root method elaborated: specificf=S_kickoff_collate leftover=1+2
//
//KiwiC: front end input processing of class or method called Testbench
//
//root_compiler: start elaborating class 'Testbench'
//
//elaborating class 'Testbench'
//
//compiling static method as entry point: style=Root idl=Testbench/Main
//
//Performing root elaboration of method Main
//
//KiwiC start_thread (or entry point) id=Main10
//
//root_compiler class done: Testbench
//
//Report of all settings used from the recipe or command line:
//
//   cil-uwind-budget=10000
//
//   kiwic-finish=enable
//
//   kiwic-cil-dump=combined
//
//   kiwic-kcode-dump=enable
//
//   array-4d-name=KIWIARRAY4D
//
//   array-3d-name=KIWIARRAY3D
//
//   array-2d-name=KIWIARRAY2D
//
//   kiwi-dll=Kiwi.dll
//
//   kiwic-dll=Kiwic.dll
//
//   kiwic-zerolength-arrays=disable
//
//   kiwic-fpgaconsole-default=enable
//
//   postgen-optimise=enable
//
//   gtrace-loglevel=20
//
//   intcil-loglevel=20
//
//   firstpass-loglevel=20
//
//   root=$attributeroot
//
//   srcfile=cuckoo_hash_demo.exe
//
//END OF KIWIC REPORT FILE
//

//----------------------------------------------------------

//Report from enumbers:::
//Concise expression alias report.
//
//  -- No expression aliases to report
//

//----------------------------------------------------------

//Report from restructure2:::
//Offchip Load/Store (and other) Ports = Nothing to Report
//

//----------------------------------------------------------

//Report from restructure2:::
//Restructure Technology Settings
//*---------------------------+---------+---------------------------------------------------------------------------------*
//| Key                       | Value   | Description                                                                     |
//*---------------------------+---------+---------------------------------------------------------------------------------*
//| int_flr_mul               | -3000   |                                                                                 |
//| fp_fl_dp_div              | 5       |                                                                                 |
//| fp_fl_dp_add              | 4       |                                                                                 |
//| fp_fl_dp_mul              | 3       |                                                                                 |
//| fp_fl_sp_div              | 5       |                                                                                 |
//| fp_fl_sp_add              | 4       |                                                                                 |
//| fp_fl_sp_mul              | 3       |                                                                                 |
//| res2-loadstore-port-count | 0       |                                                                                 |
//| max_no_fp_muls            | 6       | Maximum number of adders and subtractors (or combos) to instantiate per thread. |
//| max_no_fp_muls            | 6       | Maximum number of f/p dividers to instantiate per thread.                       |
//| max_no_int_muls           | 3       | Maximum number of int multipliers to instantiate per thread.                    |
//| max_no_fp_divs            | 2       | Maximum number of f/p dividers to instantiate per thread.                       |
//| max_no_int_divs           | 2       | Maximum number of int dividers to instantiate per thread.                       |
//| res2-offchip-threshold    | 1000000 |                                                                                 |
//| res2-combrom-threshold    | 64      |                                                                                 |
//| res2-combram-threshold    | 32      |                                                                                 |
//| res2-regfile-threshold    | 8       |                                                                                 |
//*---------------------------+---------+---------------------------------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//PC codings points for xpc10 
//*---------------------+------+--------------+------+------+-------+-----+-------------+------*
//| gb-flag/Pause       | eno  | hwm          | root | exec | start | end | antecedants | next |
//*---------------------+------+--------------+------+------+-------+-----+-------------+------*
//|   X0:"xpc10:start0" | 900  | hwm=0.0.0    | 0    | 0    | -     | -   | ---         | 1    |
//|   X1:"xpc10:1"      | 901  | hwm=0.0.0    | 1    | 1    | -     | -   | ---         | 2    |
//|   X2:"xpc10:2"      | 902  | hwm=0.0.0    | 2    | 2    | -     | -   | ---         | 3    |
//|   X3:"xpc10:3"      | 903  | hwm=0.0.0    | 3    | 3    | -     | -   | ---         | 4    |
//|   X4:"xpc10:4"      | 904  | hwm=0.0.0    | 4    | 4    | -     | -   | ---         | 5    |
//|   X5:"xpc10:5"      | 905  | hwm=0.0.0    | 5    | 5    | -     | -   | ---         | 6    |
//|   X6:"xpc10:6"      | 906  | hwm=0.0.0    | 6    | 6    | -     | -   | ---         | 7    |
//|   X7:"xpc10:7"      | 907  | hwm=0.0.0    | 7    | 7    | -     | -   | ---         | 8    |
//|   X8:"xpc10:8"      | 908  | hwm=0.0.0    | 8    | 8    | -     | -   | ---         | 9    |
//|   X9:"xpc10:9"      | 909  | hwm=0.0.0    | 9    | 9    | -     | -   | ---         | 10   |
//|   X10:"xpc10:10"    | 910  | hwm=0.0.0    | 10   | 10   | -     | -   | ---         | 11   |
//|   X11:"xpc10:11"    | 911  | hwm=0.0.0    | 11   | 11   | -     | -   | ---         | 12   |
//|   X12:"xpc10:12"    | 912  | hwm=0.0.0    | 12   | 12   | -     | -   | ---         | 13   |
//|   X13:"xpc10:13"    | 913  | hwm=0.0.0    | 13   | 13   | -     | -   | ---         | 14   |
//|   X14:"xpc10:14"    | 914  | hwm=0.0.0    | 14   | 14   | -     | -   | ---         | 15   |
//|   X15:"xpc10:15"    | 915  | hwm=0.0.0    | 15   | 15   | -     | -   | ---         | 16   |
//|   X16:"xpc10:16"    | 916  | hwm=0.0.0    | 16   | 16   | -     | -   | ---         | 17   |
//|   X17:"xpc10:17"    | 917  | hwm=0.0.0    | 17   | 17   | -     | -   | ---         | 18   |
//|   X18:"xpc10:18"    | 918  | hwm=0.0.0    | 18   | 18   | -     | -   | ---         | 19   |
//|   X19:"xpc10:19"    | 919  | hwm=0.0.0    | 19   | 19   | -     | -   | ---         | 20   |
//|   X20:"xpc10:20"    | 936  | hwm=0.0.0    | 20   | 20   | -     | -   | ---         | 65   |
//|   X20:"xpc10:20"    | 935  | hwm=0.0.1    | 20   | 20   | 36    | 36  | ---         | 549  |
//|   X20:"xpc10:20"    | 934  | hwm=0.0.1    | 20   | 20   | 35    | 35  | ---         | 547  |
//|   X20:"xpc10:20"    | 933  | hwm=0.0.1    | 20   | 20   | 34    | 34  | ---         | 544  |
//|   X20:"xpc10:20"    | 932  | hwm=0.0.1    | 20   | 20   | 33    | 33  | ---         | 540  |
//|   X20:"xpc10:20"    | 931  | hwm=0.0.1    | 20   | 20   | 32    | 32  | ---         | 571  |
//|   X20:"xpc10:20"    | 930  | hwm=0.0.1    | 20   | 20   | 31    | 31  | ---         | 565  |
//|   X20:"xpc10:20"    | 929  | hwm=0.0.1    | 20   | 20   | 30    | 30  | ---         | 558  |
//|   X20:"xpc10:20"    | 928  | hwm=0.0.1    | 20   | 20   | 29    | 29  | ---         | 550  |
//|   X20:"xpc10:20"    | 927  | hwm=0.0.1    | 20   | 20   | 28    | 28  | ---         | 609  |
//|   X20:"xpc10:20"    | 926  | hwm=0.0.1    | 20   | 20   | 27    | 27  | ---         | 599  |
//|   X20:"xpc10:20"    | 925  | hwm=0.0.1    | 20   | 20   | 26    | 26  | ---         | 588  |
//|   X20:"xpc10:20"    | 924  | hwm=0.0.1    | 20   | 20   | 25    | 25  | ---         | 576  |
//|   X20:"xpc10:20"    | 923  | hwm=0.0.1    | 20   | 20   | 24    | 24  | ---         | 37   |
//|   X20:"xpc10:20"    | 922  | hwm=0.0.1    | 20   | 20   | 23    | 23  | ---         | 37   |
//|   X20:"xpc10:20"    | 921  | hwm=0.0.1    | 20   | 20   | 22    | 22  | ---         | 37   |
//|   X20:"xpc10:20"    | 920  | hwm=0.0.1    | 20   | 20   | 21    | 21  | ---         | 37   |
//|   X21:"xpc10:21"    | 949  | hwm=0.0.0    | 37   | 37   | -     | -   | ---         | 65   |
//|   X21:"xpc10:21"    | 948  | hwm=0.0.1    | 37   | 37   | 49    | 49  | ---         | 549  |
//|   X21:"xpc10:21"    | 947  | hwm=0.0.1    | 37   | 37   | 48    | 48  | ---         | 547  |
//|   X21:"xpc10:21"    | 946  | hwm=0.0.1    | 37   | 37   | 47    | 47  | ---         | 544  |
//|   X21:"xpc10:21"    | 945  | hwm=0.0.1    | 37   | 37   | 46    | 46  | ---         | 540  |
//|   X21:"xpc10:21"    | 944  | hwm=0.0.1    | 37   | 37   | 45    | 45  | ---         | 571  |
//|   X21:"xpc10:21"    | 943  | hwm=0.0.1    | 37   | 37   | 44    | 44  | ---         | 565  |
//|   X21:"xpc10:21"    | 942  | hwm=0.0.1    | 37   | 37   | 43    | 43  | ---         | 558  |
//|   X21:"xpc10:21"    | 941  | hwm=0.0.1    | 37   | 37   | 42    | 42  | ---         | 550  |
//|   X21:"xpc10:21"    | 940  | hwm=0.0.1    | 37   | 37   | 41    | 41  | ---         | 50   |
//|   X21:"xpc10:21"    | 939  | hwm=0.0.1    | 37   | 37   | 40    | 40  | ---         | 50   |
//|   X21:"xpc10:21"    | 938  | hwm=0.0.1    | 37   | 37   | 39    | 39  | ---         | 50   |
//|   X21:"xpc10:21"    | 937  | hwm=0.0.1    | 37   | 37   | 38    | 38  | ---         | 50   |
//|   X22:"xpc10:22"    | 958  | hwm=0.0.0    | 50   | 50   | -     | -   | ---         | 65   |
//|   X22:"xpc10:22"    | 957  | hwm=0.0.1    | 50   | 50   | 58    | 58  | ---         | 549  |
//|   X22:"xpc10:22"    | 956  | hwm=0.0.1    | 50   | 50   | 57    | 57  | ---         | 547  |
//|   X22:"xpc10:22"    | 955  | hwm=0.0.1    | 50   | 50   | 56    | 56  | ---         | 544  |
//|   X22:"xpc10:22"    | 954  | hwm=0.0.1    | 50   | 50   | 55    | 55  | ---         | 540  |
//|   X22:"xpc10:22"    | 953  | hwm=0.0.1    | 50   | 50   | 54    | 54  | ---         | 59   |
//|   X22:"xpc10:22"    | 952  | hwm=0.0.1    | 50   | 50   | 53    | 53  | ---         | 59   |
//|   X22:"xpc10:22"    | 951  | hwm=0.0.1    | 50   | 50   | 52    | 52  | ---         | 59   |
//|   X22:"xpc10:22"    | 950  | hwm=0.0.1    | 50   | 50   | 51    | 51  | ---         | 59   |
//|   X23:"xpc10:23"    | 963  | hwm=0.0.0    | 59   | 59   | -     | -   | ---         | 65   |
//|   X23:"xpc10:23"    | 962  | hwm=0.0.1    | 59   | 59   | 63    | 63  | ---         | 64   |
//|   X23:"xpc10:23"    | 961  | hwm=0.0.1    | 59   | 59   | 62    | 62  | ---         | 64   |
//|   X23:"xpc10:23"    | 960  | hwm=0.0.1    | 59   | 59   | 61    | 61  | ---         | 64   |
//|   X23:"xpc10:23"    | 959  | hwm=0.0.1    | 59   | 59   | 60    | 60  | ---         | 64   |
//|   X24:"xpc10:24"    | 964  | hwm=0.0.0    | 64   | 64   | -     | -   | ---         | 65   |
//|   X25:"xpc10:25"    | 982  | hwm=0.0.1    | 65   | 65   | 81    | 81  | ---         | 539  |
//|   X25:"xpc10:25"    | 981  | hwm=0.0.1    | 65   | 65   | 80    | 80  | ---         | 537  |
//|   X25:"xpc10:25"    | 980  | hwm=0.0.1    | 65   | 65   | 79    | 79  | ---         | 534  |
//|   X25:"xpc10:25"    | 979  | hwm=0.0.1    | 65   | 65   | 78    | 78  | ---         | 528  |
//|   X25:"xpc10:25"    | 978  | hwm=0.0.1    | 65   | 65   | 77    | 77  | ---         | 539  |
//|   X25:"xpc10:25"    | 977  | hwm=0.0.1    | 65   | 65   | 76    | 76  | ---         | 537  |
//|   X25:"xpc10:25"    | 976  | hwm=0.0.1    | 65   | 65   | 75    | 75  | ---         | 534  |
//|   X25:"xpc10:25"    | 975  | hwm=0.0.1    | 65   | 65   | 74    | 74  | ---         | 528  |
//|   X25:"xpc10:25"    | 974  | hwm=0.0.1    | 65   | 65   | 73    | 73  | ---         | 539  |
//|   X25:"xpc10:25"    | 973  | hwm=0.0.1    | 65   | 65   | 72    | 72  | ---         | 537  |
//|   X25:"xpc10:25"    | 972  | hwm=0.0.1    | 65   | 65   | 71    | 71  | ---         | 534  |
//|   X25:"xpc10:25"    | 971  | hwm=0.0.1    | 65   | 65   | 70    | 70  | ---         | 528  |
//|   X25:"xpc10:25"    | 970  | hwm=0.0.1    | 65   | 65   | 69    | 69  | ---         | 539  |
//|   X25:"xpc10:25"    | 969  | hwm=0.0.1    | 65   | 65   | 68    | 68  | ---         | 537  |
//|   X25:"xpc10:25"    | 968  | hwm=0.0.1    | 65   | 65   | 67    | 67  | ---         | 534  |
//|   X25:"xpc10:25"    | 967  | hwm=0.0.1    | 65   | 65   | 66    | 66  | ---         | 528  |
//|   X25:"xpc10:25"    | 966  | hwm=0.0.0    | 65   | 65   | -     | -   | ---         | 82   |
//|   X25:"xpc10:25"    | 965  | hwm=0.0.0    | 65   | 65   | -     | -   | ---         | 65   |
//|   X26:"xpc10:26"    | 983  | hwm=0.0.0    | 82   | 82   | -     | -   | ---         | 83   |
//|   X27:"xpc10:27"    | 984  | hwm=0.0.0    | 83   | 83   | -     | -   | ---         | 84   |
//|   X28:"xpc10:28"    | 985  | hwm=0.0.0    | 84   | 84   | -     | -   | ---         | 85   |
//|   X29:"xpc10:29"    | 986  | hwm=0.0.0    | 85   | 85   | -     | -   | ---         | 86   |
//|   X30:"xpc10:30"    | 988  | hwm=0.0.0    | 86   | 86   | -     | -   | ---         | 244  |
//|   X30:"xpc10:30"    | 987  | hwm=0.0.0    | 86   | 86   | -     | -   | ---         | 87   |
//|   X31:"xpc10:31"    | 989  | hwm=0.0.0    | 87   | 87   | -     | -   | ---         | 88   |
//|   X32:"xpc10:32"    | 990  | hwm=0.0.0    | 88   | 88   | -     | -   | ---         | 89   |
//|   X33:"xpc10:33"    | 991  | hwm=0.0.0    | 89   | 89   | -     | -   | ---         | 90   |
//|   X34:"xpc10:34"    | 992  | hwm=0.0.0    | 90   | 90   | -     | -   | ---         | 91   |
//|   X35:"xpc10:35"    | 993  | hwm=0.0.0    | 91   | 91   | -     | -   | ---         | 92   |
//|   X36:"xpc10:36"    | 994  | hwm=0.0.0    | 92   | 92   | -     | -   | ---         | 93   |
//|   X37:"xpc10:37"    | 995  | hwm=0.0.0    | 93   | 93   | -     | -   | ---         | 94   |
//|   X38:"xpc10:38"    | 996  | hwm=0.0.0    | 94   | 94   | -     | -   | ---         | 95   |
//|   X39:"xpc10:39"    | 998  | hwm=0.0.0    | 95   | 95   | -     | -   | ---         | 103  |
//|   X39:"xpc10:39"    | 997  | hwm=0.0.0    | 95   | 95   | -     | -   | ---         | 96   |
//|   X40:"xpc10:40"    | 1001 | hwm=0.0.0    | 96   | 96   | -     | -   | ---         | 98   |
//|   X40:"xpc10:40"    | 1000 | hwm=0.0.0    | 96   | 96   | -     | -   | ---         | 98   |
//|   X40:"xpc10:40"    | 999  | hwm=0.0.0    | 96   | 96   | -     | -   | ---         | 97   |
//|   X41:"xpc10:41"    | 1002 | hwm=0.0.0    | 97   | 97   | -     | -   | ---         | 98   |
//|   X42:"xpc10:42"    | 1003 | hwm=0.0.0    | 98   | 98   | -     | -   | ---         | 99   |
//|   X43:"xpc10:43"    | 1005 | hwm=0.0.0    | 99   | 99   | -     | -   | ---         | 90   |
//|   X43:"xpc10:43"    | 1004 | hwm=0.0.0    | 99   | 99   | -     | -   | ---         | 100  |
//|   X44:"xpc10:44"    | 1006 | hwm=0.0.0    | 100  | 100  | -     | -   | ---         | 101  |
//|   X45:"xpc10:45"    | 1007 | hwm=0.0.0    | 101  | 101  | -     | -   | ---         | 102  |
//|   X46:"xpc10:46"    | 1008 | hwm=0.0.0    | 102  | 102  | -     | -   | ---         | 102  |
//|   X47:"xpc10:47"    | 1009 | hwm=0.0.0    | 103  | 103  | -     | -   | ---         | 104  |
//|   X48:"xpc10:48"    | 1010 | hwm=0.0.0    | 104  | 104  | -     | -   | ---         | 105  |
//|   X49:"xpc10:49"    | 1011 | hwm=0.0.0    | 105  | 105  | -     | -   | ---         | 106  |
//|   X50:"xpc10:50"    | 1013 | hwm=0.64.0   | 106  | 170  | 107   | 170 | ---         | 236  |
//|   X50:"xpc10:50"    | 1012 | hwm=0.0.0    | 106  | 106  | -     | -   | ---         | 171  |
//|   X51:"xpc10:51"    | 1014 | hwm=0.64.0   | 171  | 235  | 172   | 235 | ---         | 236  |
//|   X52:"xpc10:52"    | 1017 | hwm=1.1.0    | 236  | 237  | -     | -   | ---         | 242  |
//|   X52:"xpc10:52"    | 1016 | hwm=1.1.0    | 236  | 237  | -     | -   | ---         | 239  |
//|   X52:"xpc10:52"    | 1015 | hwm=1.1.0    | 236  | 237  | -     | -   | ---         | 238  |
//|   X53:"xpc10:53"    | 1020 | hwm=0.0.0    | 238  | 238  | -     | -   | ---         | 98   |
//|   X53:"xpc10:53"    | 1019 | hwm=0.0.0    | 238  | 238  | -     | -   | ---         | 98   |
//|   X53:"xpc10:53"    | 1018 | hwm=0.0.0    | 238  | 238  | -     | -   | ---         | 97   |
//|   X54:"xpc10:54"    | 1021 | hwm=0.1.0    | 239  | 240  | 240   | 240 | ---         | 241  |
//|   X55:"xpc10:55"    | 1022 | hwm=0.0.0    | 241  | 241  | -     | -   | ---         | 238  |
//|   X56:"xpc10:56"    | 1025 | hwm=0.0.0    | 242  | 242  | -     | -   | ---         | 105  |
//|   X56:"xpc10:56"    | 1024 | hwm=0.1.0    | 242  | 243  | 243   | 243 | ---         | 239  |
//|   X56:"xpc10:56"    | 1023 | hwm=0.0.0    | 242  | 242  | -     | -   | ---         | 238  |
//|   X57:"xpc10:57"    | 1026 | hwm=0.0.0    | 244  | 244  | -     | -   | ---         | 245  |
//|   X58:"xpc10:58"    | 1027 | hwm=0.0.0    | 245  | 245  | -     | -   | ---         | 246  |
//|   X59:"xpc10:59"    | 1028 | hwm=0.0.0    | 246  | 246  | -     | -   | ---         | 247  |
//|   X60:"xpc10:60"    | 1029 | hwm=0.0.0    | 247  | 247  | -     | -   | ---         | 248  |
//|   X61:"xpc10:61"    | 1030 | hwm=0.0.0    | 248  | 248  | -     | -   | ---         | 249  |
//|   X62:"xpc10:62"    | 1033 | hwm=0.0.0    | 249  | 249  | -     | -   | ---         | 254  |
//|   X62:"xpc10:62"    | 1032 | hwm=0.0.0    | 249  | 249  | -     | -   | ---         | 250  |
//|   X62:"xpc10:62"    | 1031 | hwm=0.0.0    | 249  | 249  | -     | -   | ---         | 250  |
//|   X63:"xpc10:63"    | 1035 | hwm=0.0.0    | 250  | 250  | -     | -   | ---         | 252  |
//|   X63:"xpc10:63"    | 1034 | hwm=0.0.0    | 250  | 250  | -     | -   | ---         | 251  |
//|   X64:"xpc10:64"    | 1036 | hwm=0.0.0    | 251  | 251  | -     | -   | ---         | 252  |
//|   X65:"xpc10:65"    | 1037 | hwm=0.0.0    | 252  | 252  | -     | -   | ---         | 253  |
//|   X66:"xpc10:66"    | 1039 | hwm=0.0.0    | 253  | 253  | -     | -   | ---         | 244  |
//|   X66:"xpc10:66"    | 1038 | hwm=0.0.0    | 253  | 253  | -     | -   | ---         | 87   |
//|   X67:"xpc10:67"    | 1040 | hwm=0.0.0    | 254  | 254  | -     | -   | ---         | 255  |
//|   X68:"xpc10:68"    | 1041 | hwm=0.0.1    | 255  | 255  | 256   | 256 | ---         | 257  |
//|   X69:"xpc10:69"    | 1042 | hwm=0.0.0    | 257  | 257  | -     | -   | ---         | 258  |
//|   X70:"xpc10:70"    | 1043 | hwm=0.0.0    | 258  | 258  | -     | -   | ---         | 259  |
//|   X71:"xpc10:71"    | 1070 | hwm=0.0.0    | 259  | 259  | -     | -   | ---         | 341  |
//|   X71:"xpc10:71"    | 1069 | hwm=0.0.0    | 259  | 259  | -     | -   | ---         | 250  |
//|   X71:"xpc10:71"    | 1068 | hwm=0.0.1    | 259  | 259  | 283   | 283 | ---         | 334  |
//|   X71:"xpc10:71"    | 1067 | hwm=0.0.1    | 259  | 259  | 282   | 282 | ---         | 334  |
//|   X71:"xpc10:71"    | 1066 | hwm=0.0.1    | 259  | 259  | 281   | 281 | ---         | 334  |
//|   X71:"xpc10:71"    | 1065 | hwm=0.0.1    | 259  | 259  | 280   | 280 | ---         | 334  |
//|   X71:"xpc10:71"    | 1064 | hwm=0.0.1    | 259  | 259  | 279   | 279 | ---         | 334  |
//|   X71:"xpc10:71"    | 1063 | hwm=0.0.1    | 259  | 259  | 278   | 278 | ---         | 340  |
//|   X71:"xpc10:71"    | 1062 | hwm=0.0.1    | 259  | 259  | 277   | 277 | ---         | 338  |
//|   X71:"xpc10:71"    | 1061 | hwm=0.0.1    | 259  | 259  | 276   | 276 | ---         | 335  |
//|   X71:"xpc10:71"    | 1060 | hwm=0.0.1    | 259  | 259  | 275   | 275 | ---         | 330  |
//|   X71:"xpc10:71"    | 1059 | hwm=0.0.1    | 259  | 259  | 274   | 274 | ---         | 334  |
//|   X71:"xpc10:71"    | 1058 | hwm=0.0.1    | 259  | 259  | 273   | 273 | ---         | 340  |
//|   X71:"xpc10:71"    | 1057 | hwm=0.0.1    | 259  | 259  | 272   | 272 | ---         | 338  |
//|   X71:"xpc10:71"    | 1056 | hwm=0.0.1    | 259  | 259  | 271   | 271 | ---         | 335  |
//|   X71:"xpc10:71"    | 1055 | hwm=0.0.1    | 259  | 259  | 270   | 270 | ---         | 330  |
//|   X71:"xpc10:71"    | 1054 | hwm=0.0.1    | 259  | 259  | 269   | 269 | ---         | 334  |
//|   X71:"xpc10:71"    | 1053 | hwm=0.0.1    | 259  | 259  | 268   | 268 | ---         | 340  |
//|   X71:"xpc10:71"    | 1052 | hwm=0.0.1    | 259  | 259  | 267   | 267 | ---         | 338  |
//|   X71:"xpc10:71"    | 1051 | hwm=0.0.1    | 259  | 259  | 266   | 266 | ---         | 335  |
//|   X71:"xpc10:71"    | 1050 | hwm=0.0.1    | 259  | 259  | 265   | 265 | ---         | 330  |
//|   X71:"xpc10:71"    | 1049 | hwm=0.0.1    | 259  | 259  | 264   | 264 | ---         | 334  |
//|   X71:"xpc10:71"    | 1048 | hwm=0.0.1    | 259  | 259  | 263   | 263 | ---         | 340  |
//|   X71:"xpc10:71"    | 1047 | hwm=0.0.1    | 259  | 259  | 262   | 262 | ---         | 338  |
//|   X71:"xpc10:71"    | 1046 | hwm=0.0.1    | 259  | 259  | 261   | 261 | ---         | 335  |
//|   X71:"xpc10:71"    | 1045 | hwm=0.0.1    | 259  | 259  | 260   | 260 | ---         | 330  |
//|   X71:"xpc10:71"    | 1044 | hwm=0.0.0    | 259  | 259  | -     | -   | ---         | 284  |
//|   X72:"xpc10:72"    | 1071 | hwm=0.0.0    | 284  | 284  | -     | -   | ---         | 285  |
//|   X73:"xpc10:73"    | 1072 | hwm=0.1.0    | 285  | 286  | 286   | 286 | ---         | 287  |
//|   X74:"xpc10:74"    | 1073 | hwm=0.1.0    | 287  | 288  | 288   | 288 | ---         | 289  |
//|   X75:"xpc10:75"    | 1098 | hwm=0.0.0    | 289  | 289  | -     | -   | ---         | 323  |
//|   X75:"xpc10:75"    | 1097 | hwm=0.0.1    | 289  | 289  | 313   | 313 | ---         | 318  |
//|   X75:"xpc10:75"    | 1096 | hwm=0.0.1    | 289  | 289  | 312   | 312 | ---         | 318  |
//|   X75:"xpc10:75"    | 1095 | hwm=0.0.1    | 289  | 289  | 311   | 311 | ---         | 318  |
//|   X75:"xpc10:75"    | 1094 | hwm=0.0.1    | 289  | 289  | 310   | 310 | ---         | 318  |
//|   X75:"xpc10:75"    | 1093 | hwm=0.0.1    | 289  | 289  | 309   | 309 | ---         | 318  |
//|   X75:"xpc10:75"    | 1092 | hwm=0.0.1    | 289  | 289  | 308   | 308 | ---         | 329  |
//|   X75:"xpc10:75"    | 1091 | hwm=0.0.1    | 289  | 289  | 307   | 307 | ---         | 327  |
//|   X75:"xpc10:75"    | 1090 | hwm=0.0.1    | 289  | 289  | 306   | 306 | ---         | 324  |
//|   X75:"xpc10:75"    | 1089 | hwm=0.0.1    | 289  | 289  | 305   | 305 | ---         | 314  |
//|   X75:"xpc10:75"    | 1088 | hwm=0.0.1    | 289  | 289  | 304   | 304 | ---         | 318  |
//|   X75:"xpc10:75"    | 1087 | hwm=0.0.1    | 289  | 289  | 303   | 303 | ---         | 329  |
//|   X75:"xpc10:75"    | 1086 | hwm=0.0.1    | 289  | 289  | 302   | 302 | ---         | 327  |
//|   X75:"xpc10:75"    | 1085 | hwm=0.0.1    | 289  | 289  | 301   | 301 | ---         | 324  |
//|   X75:"xpc10:75"    | 1084 | hwm=0.0.1    | 289  | 289  | 300   | 300 | ---         | 314  |
//|   X75:"xpc10:75"    | 1083 | hwm=0.0.1    | 289  | 289  | 299   | 299 | ---         | 318  |
//|   X75:"xpc10:75"    | 1082 | hwm=0.0.1    | 289  | 289  | 298   | 298 | ---         | 329  |
//|   X75:"xpc10:75"    | 1081 | hwm=0.0.1    | 289  | 289  | 297   | 297 | ---         | 327  |
//|   X75:"xpc10:75"    | 1080 | hwm=0.0.1    | 289  | 289  | 296   | 296 | ---         | 324  |
//|   X75:"xpc10:75"    | 1079 | hwm=0.0.1    | 289  | 289  | 295   | 295 | ---         | 314  |
//|   X75:"xpc10:75"    | 1078 | hwm=0.0.1    | 289  | 289  | 294   | 294 | ---         | 318  |
//|   X75:"xpc10:75"    | 1077 | hwm=0.0.1    | 289  | 289  | 293   | 293 | ---         | 329  |
//|   X75:"xpc10:75"    | 1076 | hwm=0.0.1    | 289  | 289  | 292   | 292 | ---         | 327  |
//|   X75:"xpc10:75"    | 1075 | hwm=0.0.1    | 289  | 289  | 291   | 291 | ---         | 324  |
//|   X75:"xpc10:75"    | 1074 | hwm=0.0.1    | 289  | 289  | 290   | 290 | ---         | 314  |
//|   X76:"xpc10:76"    | 1102 | hwm=0.0.0    | 314  | 314  | -     | -   | ---         | 323  |
//|   X76:"xpc10:76"    | 1101 | hwm=0.0.1    | 314  | 314  | 317   | 317 | ---         | 318  |
//|   X76:"xpc10:76"    | 1100 | hwm=0.0.1    | 314  | 314  | 316   | 316 | ---         | 318  |
//|   X76:"xpc10:76"    | 1099 | hwm=0.0.1    | 314  | 314  | 315   | 315 | ---         | 318  |
//|   X77:"xpc10:77"    | 1103 | hwm=0.0.0    | 318  | 318  | -     | -   | ---         | 319  |
//|   X78:"xpc10:78"    | 1104 | hwm=0.0.0    | 319  | 319  | -     | -   | ---         | 320  |
//|   X79:"xpc10:79"    | 1105 | hwm=0.0.0    | 320  | 320  | -     | -   | ---         | 321  |
//|   X80:"xpc10:80"    | 1106 | hwm=0.0.0    | 321  | 321  | -     | -   | ---         | 322  |
//|   X81:"xpc10:81"    | 1107 | hwm=0.0.0    | 322  | 322  | -     | -   | ---         | 259  |
//|   X82:"xpc10:82"    | 1108 | hwm=0.0.0    | 323  | 323  | -     | -   | ---         | 320  |
//|   X83:"xpc10:83"    | 1111 | hwm=0.0.0    | 324  | 324  | -     | -   | ---         | 323  |
//|   X83:"xpc10:83"    | 1110 | hwm=0.0.1    | 324  | 324  | 326   | 326 | ---         | 318  |
//|   X83:"xpc10:83"    | 1109 | hwm=0.0.1    | 324  | 324  | 325   | 325 | ---         | 318  |
//|   X84:"xpc10:84"    | 1113 | hwm=0.0.0    | 327  | 327  | -     | -   | ---         | 323  |
//|   X84:"xpc10:84"    | 1112 | hwm=0.0.1    | 327  | 327  | 328   | 328 | ---         | 318  |
//|   X85:"xpc10:85"    | 1114 | hwm=0.0.0    | 329  | 329  | -     | -   | ---         | 323  |
//|   X86:"xpc10:86"    | 1118 | hwm=0.0.0    | 330  | 330  | -     | -   | ---         | 250  |
//|   X86:"xpc10:86"    | 1117 | hwm=0.0.1    | 330  | 330  | 333   | 333 | ---         | 334  |
//|   X86:"xpc10:86"    | 1116 | hwm=0.0.1    | 330  | 330  | 332   | 332 | ---         | 334  |
//|   X86:"xpc10:86"    | 1115 | hwm=0.0.1    | 330  | 330  | 331   | 331 | ---         | 334  |
//|   X87:"xpc10:87"    | 1120 | hwm=0.0.0    | 334  | 334  | -     | -   | ---         | 252  |
//|   X87:"xpc10:87"    | 1119 | hwm=0.0.0    | 334  | 334  | -     | -   | ---         | 251  |
//|   X88:"xpc10:88"    | 1123 | hwm=0.0.0    | 335  | 335  | -     | -   | ---         | 250  |
//|   X88:"xpc10:88"    | 1122 | hwm=0.0.1    | 335  | 335  | 337   | 337 | ---         | 334  |
//|   X88:"xpc10:88"    | 1121 | hwm=0.0.1    | 335  | 335  | 336   | 336 | ---         | 334  |
//|   X89:"xpc10:89"    | 1125 | hwm=0.0.0    | 338  | 338  | -     | -   | ---         | 250  |
//|   X89:"xpc10:89"    | 1124 | hwm=0.0.1    | 338  | 338  | 339   | 339 | ---         | 334  |
//|   X90:"xpc10:90"    | 1126 | hwm=0.0.0    | 340  | 340  | -     | -   | ---         | 250  |
//|   X91:"xpc10:91"    | 1127 | hwm=0.0.0    | 341  | 341  | -     | -   | ---         | 342  |
//|   X92:"xpc10:92"    | 1129 | hwm=0.64.0   | 342  | 406  | 343   | 406 | ---         | 472  |
//|   X92:"xpc10:92"    | 1128 | hwm=0.0.0    | 342  | 342  | -     | -   | ---         | 407  |
//|   X93:"xpc10:93"    | 1130 | hwm=0.64.0   | 407  | 471  | 408   | 471 | ---         | 472  |
//|   X94:"xpc10:94"    | 1161 | hwm=1.1.0    | 472  | 473  | -     | -   | ---         | 503  |
//|   X94:"xpc10:94"    | 1160 | hwm=1.1.0    | 472  | 473  | -     | -   | ---         | 250  |
//|   X94:"xpc10:94"    | 1159 | hwm=1.1.1    | 472  | 473  | 501   | 501 | ---         | 334  |
//|   X94:"xpc10:94"    | 1158 | hwm=1.1.1    | 472  | 473  | 500   | 500 | ---         | 334  |
//|   X94:"xpc10:94"    | 1157 | hwm=1.1.1    | 472  | 473  | 499   | 499 | ---         | 334  |
//|   X94:"xpc10:94"    | 1156 | hwm=1.1.1    | 472  | 473  | 498   | 498 | ---         | 334  |
//|   X94:"xpc10:94"    | 1155 | hwm=1.1.0    | 472  | 473  | -     | -   | ---         | 284  |
//|   X94:"xpc10:94"    | 1154 | hwm=1.1.1    | 472  | 473  | 497   | 497 | ---         | 334  |
//|   X94:"xpc10:94"    | 1153 | hwm=1.1.1    | 472  | 473  | 496   | 496 | ---         | 340  |
//|   X94:"xpc10:94"    | 1152 | hwm=1.1.1    | 472  | 473  | 495   | 495 | ---         | 338  |
//|   X94:"xpc10:94"    | 1151 | hwm=1.1.1    | 472  | 473  | 494   | 494 | ---         | 335  |
//|   X94:"xpc10:94"    | 1150 | hwm=1.1.1    | 472  | 473  | 493   | 493 | ---         | 330  |
//|   X94:"xpc10:94"    | 1149 | hwm=1.1.1    | 472  | 473  | 492   | 492 | ---         | 502  |
//|   X94:"xpc10:94"    | 1148 | hwm=1.1.1    | 472  | 473  | 491   | 491 | ---         | 334  |
//|   X94:"xpc10:94"    | 1147 | hwm=1.1.1    | 472  | 473  | 490   | 490 | ---         | 340  |
//|   X94:"xpc10:94"    | 1146 | hwm=1.1.1    | 472  | 473  | 489   | 489 | ---         | 338  |
//|   X94:"xpc10:94"    | 1145 | hwm=1.1.1    | 472  | 473  | 488   | 488 | ---         | 335  |
//|   X94:"xpc10:94"    | 1144 | hwm=1.1.1    | 472  | 473  | 487   | 487 | ---         | 330  |
//|   X94:"xpc10:94"    | 1143 | hwm=1.1.1    | 472  | 473  | 486   | 486 | ---         | 502  |
//|   X94:"xpc10:94"    | 1142 | hwm=1.1.1    | 472  | 473  | 485   | 485 | ---         | 334  |
//|   X94:"xpc10:94"    | 1141 | hwm=1.1.1    | 472  | 473  | 484   | 484 | ---         | 340  |
//|   X94:"xpc10:94"    | 1140 | hwm=1.1.1    | 472  | 473  | 483   | 483 | ---         | 338  |
//|   X94:"xpc10:94"    | 1139 | hwm=1.1.1    | 472  | 473  | 482   | 482 | ---         | 335  |
//|   X94:"xpc10:94"    | 1138 | hwm=1.1.1    | 472  | 473  | 481   | 481 | ---         | 330  |
//|   X94:"xpc10:94"    | 1137 | hwm=1.1.1    | 472  | 473  | 480   | 480 | ---         | 502  |
//|   X94:"xpc10:94"    | 1136 | hwm=1.1.1    | 472  | 473  | 479   | 479 | ---         | 334  |
//|   X94:"xpc10:94"    | 1135 | hwm=1.1.1    | 472  | 473  | 478   | 478 | ---         | 340  |
//|   X94:"xpc10:94"    | 1134 | hwm=1.1.1    | 472  | 473  | 477   | 477 | ---         | 338  |
//|   X94:"xpc10:94"    | 1133 | hwm=1.1.1    | 472  | 473  | 476   | 476 | ---         | 335  |
//|   X94:"xpc10:94"    | 1132 | hwm=1.1.1    | 472  | 473  | 475   | 475 | ---         | 330  |
//|   X94:"xpc10:94"    | 1131 | hwm=1.1.1    | 472  | 473  | 474   | 474 | ---         | 502  |
//|   X95:"xpc10:95"    | 1162 | hwm=0.0.0    | 502  | 502  | -     | -   | ---         | 284  |
//|   X96:"xpc10:96"    | 1189 | hwm=0.0.0    | 503  | 503  | -     | -   | ---         | 341  |
//|   X96:"xpc10:96"    | 1188 | hwm=0.0.0    | 503  | 503  | -     | -   | ---         | 250  |
//|   X96:"xpc10:96"    | 1187 | hwm=0.0.1    | 503  | 503  | 527   | 527 | ---         | 334  |
//|   X96:"xpc10:96"    | 1186 | hwm=0.0.1    | 503  | 503  | 526   | 526 | ---         | 334  |
//|   X96:"xpc10:96"    | 1185 | hwm=0.0.1    | 503  | 503  | 525   | 525 | ---         | 334  |
//|   X96:"xpc10:96"    | 1184 | hwm=0.0.1    | 503  | 503  | 524   | 524 | ---         | 334  |
//|   X96:"xpc10:96"    | 1183 | hwm=0.0.1    | 503  | 503  | 523   | 523 | ---         | 334  |
//|   X96:"xpc10:96"    | 1182 | hwm=0.0.1    | 503  | 503  | 522   | 522 | ---         | 340  |
//|   X96:"xpc10:96"    | 1181 | hwm=0.0.1    | 503  | 503  | 521   | 521 | ---         | 338  |
//|   X96:"xpc10:96"    | 1180 | hwm=0.0.1    | 503  | 503  | 520   | 520 | ---         | 335  |
//|   X96:"xpc10:96"    | 1179 | hwm=0.0.1    | 503  | 503  | 519   | 519 | ---         | 330  |
//|   X96:"xpc10:96"    | 1178 | hwm=0.0.1    | 503  | 503  | 518   | 518 | ---         | 334  |
//|   X96:"xpc10:96"    | 1177 | hwm=0.0.1    | 503  | 503  | 517   | 517 | ---         | 340  |
//|   X96:"xpc10:96"    | 1176 | hwm=0.0.1    | 503  | 503  | 516   | 516 | ---         | 338  |
//|   X96:"xpc10:96"    | 1175 | hwm=0.0.1    | 503  | 503  | 515   | 515 | ---         | 335  |
//|   X96:"xpc10:96"    | 1174 | hwm=0.0.1    | 503  | 503  | 514   | 514 | ---         | 330  |
//|   X96:"xpc10:96"    | 1173 | hwm=0.0.1    | 503  | 503  | 513   | 513 | ---         | 334  |
//|   X96:"xpc10:96"    | 1172 | hwm=0.0.1    | 503  | 503  | 512   | 512 | ---         | 340  |
//|   X96:"xpc10:96"    | 1171 | hwm=0.0.1    | 503  | 503  | 511   | 511 | ---         | 338  |
//|   X96:"xpc10:96"    | 1170 | hwm=0.0.1    | 503  | 503  | 510   | 510 | ---         | 335  |
//|   X96:"xpc10:96"    | 1169 | hwm=0.0.1    | 503  | 503  | 509   | 509 | ---         | 330  |
//|   X96:"xpc10:96"    | 1168 | hwm=0.0.1    | 503  | 503  | 508   | 508 | ---         | 334  |
//|   X96:"xpc10:96"    | 1167 | hwm=0.0.1    | 503  | 503  | 507   | 507 | ---         | 340  |
//|   X96:"xpc10:96"    | 1166 | hwm=0.0.1    | 503  | 503  | 506   | 506 | ---         | 338  |
//|   X96:"xpc10:96"    | 1165 | hwm=0.0.1    | 503  | 503  | 505   | 505 | ---         | 335  |
//|   X96:"xpc10:96"    | 1164 | hwm=0.0.1    | 503  | 503  | 504   | 504 | ---         | 330  |
//|   X96:"xpc10:96"    | 1163 | hwm=0.0.0    | 503  | 503  | -     | -   | ---         | 284  |
//|   X97:"xpc10:97"    | 1193 | hwm=0.0.0    | 528  | 528  | -     | -   | ---         | 532  |
//|   X97:"xpc10:97"    | 1192 | hwm=0.0.1    | 528  | 528  | 531   | 531 | ---         | 532  |
//|   X97:"xpc10:97"    | 1191 | hwm=0.0.1    | 528  | 528  | 530   | 530 | ---         | 532  |
//|   X97:"xpc10:97"    | 1190 | hwm=0.0.1    | 528  | 528  | 529   | 529 | ---         | 532  |
//|   X98:"xpc10:98"    | 1195 | hwm=0.0.0    | 532  | 532  | -     | -   | ---         | 65   |
//|   X98:"xpc10:98"    | 1194 | hwm=0.0.1    | 532  | 532  | 533   | 533 | ---         | 532  |
//|   X99:"xpc10:99"    | 1198 | hwm=0.0.0    | 534  | 534  | -     | -   | ---         | 532  |
//|   X99:"xpc10:99"    | 1197 | hwm=0.0.1    | 534  | 534  | 536   | 536 | ---         | 532  |
//|   X99:"xpc10:99"    | 1196 | hwm=0.0.1    | 534  | 534  | 535   | 535 | ---         | 532  |
//|   X100:"xpc10:100"  | 1200 | hwm=0.0.0    | 537  | 537  | -     | -   | ---         | 532  |
//|   X100:"xpc10:100"  | 1199 | hwm=0.0.1    | 537  | 537  | 538   | 538 | ---         | 532  |
//|   X101:"xpc10:101"  | 1201 | hwm=0.0.0    | 539  | 539  | -     | -   | ---         | 532  |
//|   X102:"xpc10:102"  | 1205 | hwm=0.0.0    | 540  | 540  | -     | -   | ---         | 65   |
//|   X102:"xpc10:102"  | 1204 | hwm=0.0.1    | 540  | 540  | 543   | 543 | ---         | 64   |
//|   X102:"xpc10:102"  | 1203 | hwm=0.0.1    | 540  | 540  | 542   | 542 | ---         | 64   |
//|   X102:"xpc10:102"  | 1202 | hwm=0.0.1    | 540  | 540  | 541   | 541 | ---         | 64   |
//|   X103:"xpc10:103"  | 1208 | hwm=0.0.0    | 544  | 544  | -     | -   | ---         | 65   |
//|   X103:"xpc10:103"  | 1207 | hwm=0.0.1    | 544  | 544  | 546   | 546 | ---         | 64   |
//|   X103:"xpc10:103"  | 1206 | hwm=0.0.1    | 544  | 544  | 545   | 545 | ---         | 64   |
//|   X104:"xpc10:104"  | 1210 | hwm=0.0.0    | 547  | 547  | -     | -   | ---         | 65   |
//|   X104:"xpc10:104"  | 1209 | hwm=0.0.1    | 547  | 547  | 548   | 548 | ---         | 64   |
//|   X105:"xpc10:105"  | 1211 | hwm=0.0.0    | 549  | 549  | -     | -   | ---         | 65   |
//|   X106:"xpc10:106"  | 1219 | hwm=0.0.0    | 550  | 550  | -     | -   | ---         | 65   |
//|   X106:"xpc10:106"  | 1218 | hwm=0.0.1    | 550  | 550  | 557   | 557 | ---         | 549  |
//|   X106:"xpc10:106"  | 1217 | hwm=0.0.1    | 550  | 550  | 556   | 556 | ---         | 547  |
//|   X106:"xpc10:106"  | 1216 | hwm=0.0.1    | 550  | 550  | 555   | 555 | ---         | 544  |
//|   X106:"xpc10:106"  | 1215 | hwm=0.0.1    | 550  | 550  | 554   | 554 | ---         | 540  |
//|   X106:"xpc10:106"  | 1214 | hwm=0.0.1    | 550  | 550  | 553   | 553 | ---         | 59   |
//|   X106:"xpc10:106"  | 1213 | hwm=0.0.1    | 550  | 550  | 552   | 552 | ---         | 59   |
//|   X106:"xpc10:106"  | 1212 | hwm=0.0.1    | 550  | 550  | 551   | 551 | ---         | 59   |
//|   X107:"xpc10:107"  | 1226 | hwm=0.0.0    | 558  | 558  | -     | -   | ---         | 65   |
//|   X107:"xpc10:107"  | 1225 | hwm=0.0.1    | 558  | 558  | 564   | 564 | ---         | 549  |
//|   X107:"xpc10:107"  | 1224 | hwm=0.0.1    | 558  | 558  | 563   | 563 | ---         | 547  |
//|   X107:"xpc10:107"  | 1223 | hwm=0.0.1    | 558  | 558  | 562   | 562 | ---         | 544  |
//|   X107:"xpc10:107"  | 1222 | hwm=0.0.1    | 558  | 558  | 561   | 561 | ---         | 540  |
//|   X107:"xpc10:107"  | 1221 | hwm=0.0.1    | 558  | 558  | 560   | 560 | ---         | 59   |
//|   X107:"xpc10:107"  | 1220 | hwm=0.0.1    | 558  | 558  | 559   | 559 | ---         | 59   |
//|   X108:"xpc10:108"  | 1232 | hwm=0.0.0    | 565  | 565  | -     | -   | ---         | 65   |
//|   X108:"xpc10:108"  | 1231 | hwm=0.0.1    | 565  | 565  | 570   | 570 | ---         | 549  |
//|   X108:"xpc10:108"  | 1230 | hwm=0.0.1    | 565  | 565  | 569   | 569 | ---         | 547  |
//|   X108:"xpc10:108"  | 1229 | hwm=0.0.1    | 565  | 565  | 568   | 568 | ---         | 544  |
//|   X108:"xpc10:108"  | 1228 | hwm=0.0.1    | 565  | 565  | 567   | 567 | ---         | 540  |
//|   X108:"xpc10:108"  | 1227 | hwm=0.0.1    | 565  | 565  | 566   | 566 | ---         | 59   |
//|   X109:"xpc10:109"  | 1237 | hwm=0.0.0    | 571  | 571  | -     | -   | ---         | 65   |
//|   X109:"xpc10:109"  | 1236 | hwm=0.0.1    | 571  | 571  | 575   | 575 | ---         | 549  |
//|   X109:"xpc10:109"  | 1235 | hwm=0.0.1    | 571  | 571  | 574   | 574 | ---         | 547  |
//|   X109:"xpc10:109"  | 1234 | hwm=0.0.1    | 571  | 571  | 573   | 573 | ---         | 544  |
//|   X109:"xpc10:109"  | 1233 | hwm=0.0.1    | 571  | 571  | 572   | 572 | ---         | 540  |
//|   X110:"xpc10:110"  | 1249 | hwm=0.0.0    | 576  | 576  | -     | -   | ---         | 65   |
//|   X110:"xpc10:110"  | 1248 | hwm=0.0.1    | 576  | 576  | 587   | 587 | ---         | 549  |
//|   X110:"xpc10:110"  | 1247 | hwm=0.0.1    | 576  | 576  | 586   | 586 | ---         | 547  |
//|   X110:"xpc10:110"  | 1246 | hwm=0.0.1    | 576  | 576  | 585   | 585 | ---         | 544  |
//|   X110:"xpc10:110"  | 1245 | hwm=0.0.1    | 576  | 576  | 584   | 584 | ---         | 540  |
//|   X110:"xpc10:110"  | 1244 | hwm=0.0.1    | 576  | 576  | 583   | 583 | ---         | 571  |
//|   X110:"xpc10:110"  | 1243 | hwm=0.0.1    | 576  | 576  | 582   | 582 | ---         | 565  |
//|   X110:"xpc10:110"  | 1242 | hwm=0.0.1    | 576  | 576  | 581   | 581 | ---         | 558  |
//|   X110:"xpc10:110"  | 1241 | hwm=0.0.1    | 576  | 576  | 580   | 580 | ---         | 550  |
//|   X110:"xpc10:110"  | 1240 | hwm=0.0.1    | 576  | 576  | 579   | 579 | ---         | 50   |
//|   X110:"xpc10:110"  | 1239 | hwm=0.0.1    | 576  | 576  | 578   | 578 | ---         | 50   |
//|   X110:"xpc10:110"  | 1238 | hwm=0.0.1    | 576  | 576  | 577   | 577 | ---         | 50   |
//|   X111:"xpc10:111"  | 1260 | hwm=0.0.0    | 588  | 588  | -     | -   | ---         | 65   |
//|   X111:"xpc10:111"  | 1259 | hwm=0.0.1    | 588  | 588  | 598   | 598 | ---         | 549  |
//|   X111:"xpc10:111"  | 1258 | hwm=0.0.1    | 588  | 588  | 597   | 597 | ---         | 547  |
//|   X111:"xpc10:111"  | 1257 | hwm=0.0.1    | 588  | 588  | 596   | 596 | ---         | 544  |
//|   X111:"xpc10:111"  | 1256 | hwm=0.0.1    | 588  | 588  | 595   | 595 | ---         | 540  |
//|   X111:"xpc10:111"  | 1255 | hwm=0.0.1    | 588  | 588  | 594   | 594 | ---         | 571  |
//|   X111:"xpc10:111"  | 1254 | hwm=0.0.1    | 588  | 588  | 593   | 593 | ---         | 565  |
//|   X111:"xpc10:111"  | 1253 | hwm=0.0.1    | 588  | 588  | 592   | 592 | ---         | 558  |
//|   X111:"xpc10:111"  | 1252 | hwm=0.0.1    | 588  | 588  | 591   | 591 | ---         | 550  |
//|   X111:"xpc10:111"  | 1251 | hwm=0.0.1    | 588  | 588  | 590   | 590 | ---         | 50   |
//|   X111:"xpc10:111"  | 1250 | hwm=0.0.1    | 588  | 588  | 589   | 589 | ---         | 50   |
//|   X112:"xpc10:112"  | 1270 | hwm=0.0.0    | 599  | 599  | -     | -   | ---         | 65   |
//|   X112:"xpc10:112"  | 1269 | hwm=0.0.1    | 599  | 599  | 608   | 608 | ---         | 549  |
//|   X112:"xpc10:112"  | 1268 | hwm=0.0.1    | 599  | 599  | 607   | 607 | ---         | 547  |
//|   X112:"xpc10:112"  | 1267 | hwm=0.0.1    | 599  | 599  | 606   | 606 | ---         | 544  |
//|   X112:"xpc10:112"  | 1266 | hwm=0.0.1    | 599  | 599  | 605   | 605 | ---         | 540  |
//|   X112:"xpc10:112"  | 1265 | hwm=0.0.1    | 599  | 599  | 604   | 604 | ---         | 571  |
//|   X112:"xpc10:112"  | 1264 | hwm=0.0.1    | 599  | 599  | 603   | 603 | ---         | 565  |
//|   X112:"xpc10:112"  | 1263 | hwm=0.0.1    | 599  | 599  | 602   | 602 | ---         | 558  |
//|   X112:"xpc10:112"  | 1262 | hwm=0.0.1    | 599  | 599  | 601   | 601 | ---         | 550  |
//|   X112:"xpc10:112"  | 1261 | hwm=0.0.1    | 599  | 599  | 600   | 600 | ---         | 50   |
//|   X113:"xpc10:113"  | 1279 | hwm=0.0.0    | 609  | 609  | -     | -   | ---         | 65   |
//|   X113:"xpc10:113"  | 1278 | hwm=0.0.1    | 609  | 609  | 617   | 617 | ---         | 549  |
//|   X113:"xpc10:113"  | 1277 | hwm=0.0.1    | 609  | 609  | 616   | 616 | ---         | 547  |
//|   X113:"xpc10:113"  | 1276 | hwm=0.0.1    | 609  | 609  | 615   | 615 | ---         | 544  |
//|   X113:"xpc10:113"  | 1275 | hwm=0.0.1    | 609  | 609  | 614   | 614 | ---         | 540  |
//|   X113:"xpc10:113"  | 1274 | hwm=0.0.1    | 609  | 609  | 613   | 613 | ---         | 571  |
//|   X113:"xpc10:113"  | 1273 | hwm=0.0.1    | 609  | 609  | 612   | 612 | ---         | 565  |
//|   X113:"xpc10:113"  | 1272 | hwm=0.0.1    | 609  | 609  | 611   | 611 | ---         | 558  |
//|   X113:"xpc10:113"  | 1271 | hwm=0.0.1    | 609  | 609  | 610   | 610 | ---         | 550  |
//*---------------------+------+--------------+------+------+-------+-----+-------------+------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X0:"xpc10:start0" 900 :  major_start_pcl=0   edge_private_start/end=-1/-1 exec=0 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X0:"xpc10:start0"
//res2: Thread=xpc10 state=X0:"xpc10:start0"
//*-----+-----+---------+------*
//| pc  | eno | Phaser  | Work |
//*-----+-----+---------+------*
//| 0   | -   | R0 CTRL |      |
//| 0   | 900 | R0 DATA |      |
//| 0+E | 900 | W0 DATA |      |
//*-----+-----+---------+------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X1:"xpc10:1" 901 :  major_start_pcl=1   edge_private_start/end=-1/-1 exec=1 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X1:"xpc10:1"
//res2: Thread=xpc10 state=X1:"xpc10:1"
//*-----+-----+---------+-----------------------------------------*
//| pc  | eno | Phaser  | Work                                    |
//*-----+-----+---------+-----------------------------------------*
//| 1   | -   | R0 CTRL |                                         |
//| 1   | 901 | R0 DATA |                                         |
//| 1+E | 901 | W0 DATA |  PLI:Cuckoo cache testben...  W/P:Start |
//*-----+-----+---------+-----------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X2:"xpc10:2" 902 :  major_start_pcl=2   edge_private_start/end=-1/-1 exec=2 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X2:"xpc10:2"
//res2: Thread=xpc10 state=X2:"xpc10:2"
//*-----+-----+---------+------*
//| pc  | eno | Phaser  | Work |
//*-----+-----+---------+------*
//| 2   | -   | R0 CTRL |      |
//| 2   | 902 | R0 DATA |      |
//| 2+E | 902 | W0 DATA |      |
//*-----+-----+---------+------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X3:"xpc10:3" 903 :  major_start_pcl=3   edge_private_start/end=-1/-1 exec=3 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X3:"xpc10:3"
//res2: Thread=xpc10 state=X3:"xpc10:3"
//*-----+-----+---------+------*
//| pc  | eno | Phaser  | Work |
//*-----+-----+---------+------*
//| 3   | -   | R0 CTRL |      |
//| 3   | 903 | R0 DATA |      |
//| 3+E | 903 | W0 DATA |      |
//*-----+-----+---------+------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X4:"xpc10:4" 904 :  major_start_pcl=4   edge_private_start/end=-1/-1 exec=4 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X4:"xpc10:4"
//res2: Thread=xpc10 state=X4:"xpc10:4"
//*-----+-----+---------+----------------------------------------------------*
//| pc  | eno | Phaser  | Work                                               |
//*-----+-----+---------+----------------------------------------------------*
//| 4   | -   | R0 CTRL |                                                    |
//| 4   | 904 | R0 DATA |                                                    |
//| 4+E | 904 | W0 DATA | @_SINT/CC/SCALbx24_waycap te=te:4 scalarw(S'8192I) |
//*-----+-----+---------+----------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X5:"xpc10:5" 905 :  major_start_pcl=5   edge_private_start/end=-1/-1 exec=5 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X5:"xpc10:5"
//res2: Thread=xpc10 state=X5:"xpc10:5"
//*-----+-----+---------+------*
//| pc  | eno | Phaser  | Work |
//*-----+-----+---------+------*
//| 5   | -   | R0 CTRL |      |
//| 5   | 905 | R0 DATA |      |
//| 5+E | 905 | W0 DATA |      |
//*-----+-----+---------+------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X6:"xpc10:6" 906 :  major_start_pcl=6   edge_private_start/end=-1/-1 exec=6 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X6:"xpc10:6"
//res2: Thread=xpc10 state=X6:"xpc10:6"
//*-----+-----+---------+------*
//| pc  | eno | Phaser  | Work |
//*-----+-----+---------+------*
//| 6   | -   | R0 CTRL |      |
//| 6   | 906 | R0 DATA |      |
//| 6+E | 906 | W0 DATA |      |
//*-----+-----+---------+------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X7:"xpc10:7" 907 :  major_start_pcl=7   edge_private_start/end=-1/-1 exec=7 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X7:"xpc10:7"
//res2: Thread=xpc10 state=X7:"xpc10:7"
//*-----+-----+---------+------*
//| pc  | eno | Phaser  | Work |
//*-----+-----+---------+------*
//| 7   | -   | R0 CTRL |      |
//| 7   | 907 | R0 DATA |      |
//| 7+E | 907 | W0 DATA |      |
//*-----+-----+---------+------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X8:"xpc10:8" 908 :  major_start_pcl=8   edge_private_start/end=-1/-1 exec=8 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X8:"xpc10:8"
//res2: Thread=xpc10 state=X8:"xpc10:8"
//*-----+-----+---------+------*
//| pc  | eno | Phaser  | Work |
//*-----+-----+---------+------*
//| 8   | -   | R0 CTRL |      |
//| 8   | 908 | R0 DATA |      |
//| 8+E | 908 | W0 DATA |      |
//*-----+-----+---------+------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X9:"xpc10:9" 909 :  major_start_pcl=9   edge_private_start/end=-1/-1 exec=9 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X9:"xpc10:9"
//res2: Thread=xpc10 state=X9:"xpc10:9"
//*-----+-----+---------+------*
//| pc  | eno | Phaser  | Work |
//*-----+-----+---------+------*
//| 9   | -   | R0 CTRL |      |
//| 9   | 909 | R0 DATA |      |
//| 9+E | 909 | W0 DATA |      |
//*-----+-----+---------+------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X10:"xpc10:10" 910 :  major_start_pcl=10   edge_private_start/end=-1/-1 exec=10 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X10:"xpc10:10"
//res2: Thread=xpc10 state=X10:"xpc10:10"
//*------+-----+---------+------*
//| pc   | eno | Phaser  | Work |
//*------+-----+---------+------*
//| 10   | -   | R0 CTRL |      |
//| 10   | 910 | R0 DATA |      |
//| 10+E | 910 | W0 DATA |      |
//*------+-----+---------+------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X11:"xpc10:11" 911 :  major_start_pcl=11   edge_private_start/end=-1/-1 exec=11 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X11:"xpc10:11"
//res2: Thread=xpc10 state=X11:"xpc10:11"
//*------+-----+---------+------*
//| pc   | eno | Phaser  | Work |
//*------+-----+---------+------*
//| 11   | -   | R0 CTRL |      |
//| 11   | 911 | R0 DATA |      |
//| 11+E | 911 | W0 DATA |      |
//*------+-----+---------+------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X12:"xpc10:12" 912 :  major_start_pcl=12   edge_private_start/end=-1/-1 exec=12 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X12:"xpc10:12"
//res2: Thread=xpc10 state=X12:"xpc10:12"
//*------+-----+---------+------*
//| pc   | eno | Phaser  | Work |
//*------+-----+---------+------*
//| 12   | -   | R0 CTRL |      |
//| 12   | 912 | R0 DATA |      |
//| 12+E | 912 | W0 DATA |      |
//*------+-----+---------+------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X13:"xpc10:13" 913 :  major_start_pcl=13   edge_private_start/end=-1/-1 exec=13 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X13:"xpc10:13"
//res2: Thread=xpc10 state=X13:"xpc10:13"
//*------+-----+---------+------*
//| pc   | eno | Phaser  | Work |
//*------+-----+---------+------*
//| 13   | -   | R0 CTRL |      |
//| 13   | 913 | R0 DATA |      |
//| 13+E | 913 | W0 DATA |      |
//*------+-----+---------+------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X14:"xpc10:14" 914 :  major_start_pcl=14   edge_private_start/end=-1/-1 exec=14 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X14:"xpc10:14"
//res2: Thread=xpc10 state=X14:"xpc10:14"
//*------+-----+---------+------*
//| pc   | eno | Phaser  | Work |
//*------+-----+---------+------*
//| 14   | -   | R0 CTRL |      |
//| 14   | 914 | R0 DATA |      |
//| 14+E | 914 | W0 DATA |      |
//*------+-----+---------+------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X15:"xpc10:15" 915 :  major_start_pcl=15   edge_private_start/end=-1/-1 exec=15 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X15:"xpc10:15"
//res2: Thread=xpc10 state=X15:"xpc10:15"
//*------+-----+---------+------*
//| pc   | eno | Phaser  | Work |
//*------+-----+---------+------*
//| 15   | -   | R0 CTRL |      |
//| 15   | 915 | R0 DATA |      |
//| 15+E | 915 | W0 DATA |      |
//*------+-----+---------+------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X16:"xpc10:16" 916 :  major_start_pcl=16   edge_private_start/end=-1/-1 exec=16 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X16:"xpc10:16"
//res2: Thread=xpc10 state=X16:"xpc10:16"
//*------+-----+---------+------*
//| pc   | eno | Phaser  | Work |
//*------+-----+---------+------*
//| 16   | -   | R0 CTRL |      |
//| 16   | 916 | R0 DATA |      |
//| 16+E | 916 | W0 DATA |      |
//*------+-----+---------+------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X17:"xpc10:17" 917 :  major_start_pcl=17   edge_private_start/end=-1/-1 exec=17 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X17:"xpc10:17"
//res2: Thread=xpc10 state=X17:"xpc10:17"
//*------+-----+---------+------*
//| pc   | eno | Phaser  | Work |
//*------+-----+---------+------*
//| 17   | -   | R0 CTRL |      |
//| 17   | 917 | R0 DATA |      |
//| 17+E | 917 | W0 DATA |      |
//*------+-----+---------+------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X18:"xpc10:18" 918 :  major_start_pcl=18   edge_private_start/end=-1/-1 exec=18 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X18:"xpc10:18"
//res2: Thread=xpc10 state=X18:"xpc10:18"
//*------+-----+---------+------*
//| pc   | eno | Phaser  | Work |
//*------+-----+---------+------*
//| 18   | -   | R0 CTRL |      |
//| 18   | 918 | R0 DATA |      |
//| 18+E | 918 | W0 DATA |      |
//*------+-----+---------+------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X19:"xpc10:19" 919 :  major_start_pcl=19   edge_private_start/end=-1/-1 exec=19 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X19:"xpc10:19"
//res2: Thread=xpc10 state=X19:"xpc10:19"
//*------+-----+---------+-------------------------------------------------------------------*
//| pc   | eno | Phaser  | Work                                                              |
//*------+-----+---------+-------------------------------------------------------------------*
//| 19   | -   | R0 CTRL |                                                                   |
//| 19   | 919 | R0 DATA |                                                                   |
//| 19+E | 919 | W0 DATA | TCCl0.12_V_1 te=te:19 scalarw(0) TCCl0.12_V_0 te=te:19 scalarw(0) |
//*------+-----+---------+-------------------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X20:"xpc10:20" 936 :  major_start_pcl=20   edge_private_start/end=-1/-1 exec=20 (dend=0)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X20:"xpc10:20" 935 :  major_start_pcl=20   edge_private_start/end=36/36 exec=20 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X20:"xpc10:20" 934 :  major_start_pcl=20   edge_private_start/end=35/35 exec=20 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X20:"xpc10:20" 933 :  major_start_pcl=20   edge_private_start/end=34/34 exec=20 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X20:"xpc10:20" 932 :  major_start_pcl=20   edge_private_start/end=33/33 exec=20 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X20:"xpc10:20" 931 :  major_start_pcl=20   edge_private_start/end=32/32 exec=20 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X20:"xpc10:20" 930 :  major_start_pcl=20   edge_private_start/end=31/31 exec=20 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X20:"xpc10:20" 929 :  major_start_pcl=20   edge_private_start/end=30/30 exec=20 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X20:"xpc10:20" 928 :  major_start_pcl=20   edge_private_start/end=29/29 exec=20 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X20:"xpc10:20" 927 :  major_start_pcl=20   edge_private_start/end=28/28 exec=20 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X20:"xpc10:20" 926 :  major_start_pcl=20   edge_private_start/end=27/27 exec=20 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X20:"xpc10:20" 925 :  major_start_pcl=20   edge_private_start/end=26/26 exec=20 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X20:"xpc10:20" 924 :  major_start_pcl=20   edge_private_start/end=25/25 exec=20 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X20:"xpc10:20" 923 :  major_start_pcl=20   edge_private_start/end=24/24 exec=20 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X20:"xpc10:20" 922 :  major_start_pcl=20   edge_private_start/end=23/23 exec=20 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X20:"xpc10:20" 921 :  major_start_pcl=20   edge_private_start/end=22/22 exec=20 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X20:"xpc10:20" 920 :  major_start_pcl=20   edge_private_start/end=21/21 exec=20 (dend=1)
//Simple greedy schedule for res2: Thread=xpc10 state=X20:"xpc10:20"
//res2: Thread=xpc10 state=X20:"xpc10:20"
//*------+-----+---------+----------------------------------------------------------------------------------*
//| pc   | eno | Phaser  | Work                                                                             |
//*------+-----+---------+----------------------------------------------------------------------------------*
//| 20   | -   | R0 CTRL |                                                                                  |
//| 20   | 920 | R0 DATA |                                                                                  |
//| 20+E | 920 | W0 DATA | TCCl0.12_V_1 te=te:20 scalarw(1) @_SINT/CC/MAPR10NoCE3_ARA0 te=te:20 write(0, 0) |
//| 21   | 920 | W1 DATA |                                                                                  |
//| 20   | 921 | R0 DATA |                                                                                  |
//| 20+E | 921 | W0 DATA | TCCl0.12_V_1 te=te:20 scalarw(1) @_SINT/CC/MAPR10NoCE2_ARA0 te=te:20 write(0, 0) |
//| 22   | 921 | W1 DATA |                                                                                  |
//| 20   | 922 | R0 DATA |                                                                                  |
//| 20+E | 922 | W0 DATA | TCCl0.12_V_1 te=te:20 scalarw(1) @_SINT/CC/MAPR10NoCE1_ARA0 te=te:20 write(0, 0) |
//| 23   | 922 | W1 DATA |                                                                                  |
//| 20   | 923 | R0 DATA |                                                                                  |
//| 20+E | 923 | W0 DATA | TCCl0.12_V_1 te=te:20 scalarw(1) @_SINT/CC/MAPR10NoCE0_ARA0 te=te:20 write(0, 0) |
//| 24   | 923 | W1 DATA |                                                                                  |
//| 20   | 924 | R0 DATA |                                                                                  |
//| 20+E | 924 | W0 DATA | TCCl0.12_V_1 te=te:20 scalarw(1) @_SINT/CC/MAPR10NoCE3_ARA0 te=te:20 write(0, 0) |
//| 25   | 924 | W1 DATA |                                                                                  |
//| 20   | 925 | R0 DATA |                                                                                  |
//| 20+E | 925 | W0 DATA | TCCl0.12_V_1 te=te:20 scalarw(1) @_SINT/CC/MAPR10NoCE2_ARA0 te=te:20 write(0, 0) |
//| 26   | 925 | W1 DATA |                                                                                  |
//| 20   | 926 | R0 DATA |                                                                                  |
//| 20+E | 926 | W0 DATA | TCCl0.12_V_1 te=te:20 scalarw(1) @_SINT/CC/MAPR10NoCE1_ARA0 te=te:20 write(0, 0) |
//| 27   | 926 | W1 DATA |                                                                                  |
//| 20   | 927 | R0 DATA |                                                                                  |
//| 20+E | 927 | W0 DATA | TCCl0.12_V_1 te=te:20 scalarw(1) @_SINT/CC/MAPR10NoCE0_ARA0 te=te:20 write(0, 0) |
//| 28   | 927 | W1 DATA |                                                                                  |
//| 20   | 928 | R0 DATA |                                                                                  |
//| 20+E | 928 | W0 DATA | TCCl0.12_V_1 te=te:20 scalarw(2) @_SINT/CC/MAPR10NoCE3_ARA0 te=te:20 write(0, 0) |
//| 29   | 928 | W1 DATA |                                                                                  |
//| 20   | 929 | R0 DATA |                                                                                  |
//| 20+E | 929 | W0 DATA | TCCl0.12_V_1 te=te:20 scalarw(2) @_SINT/CC/MAPR10NoCE2_ARA0 te=te:20 write(0, 0) |
//| 30   | 929 | W1 DATA |                                                                                  |
//| 20   | 930 | R0 DATA |                                                                                  |
//| 20+E | 930 | W0 DATA | TCCl0.12_V_1 te=te:20 scalarw(2) @_SINT/CC/MAPR10NoCE1_ARA0 te=te:20 write(0, 0) |
//| 31   | 930 | W1 DATA |                                                                                  |
//| 20   | 931 | R0 DATA |                                                                                  |
//| 20+E | 931 | W0 DATA | TCCl0.12_V_1 te=te:20 scalarw(2) @_SINT/CC/MAPR10NoCE0_ARA0 te=te:20 write(0, 0) |
//| 32   | 931 | W1 DATA |                                                                                  |
//| 20   | 932 | R0 DATA |                                                                                  |
//| 20+E | 932 | W0 DATA | TCCl0.12_V_1 te=te:20 scalarw(3) @_SINT/CC/MAPR10NoCE3_ARA0 te=te:20 write(0, 0) |
//| 33   | 932 | W1 DATA |                                                                                  |
//| 20   | 933 | R0 DATA |                                                                                  |
//| 20+E | 933 | W0 DATA | TCCl0.12_V_1 te=te:20 scalarw(3) @_SINT/CC/MAPR10NoCE2_ARA0 te=te:20 write(0, 0) |
//| 34   | 933 | W1 DATA |                                                                                  |
//| 20   | 934 | R0 DATA |                                                                                  |
//| 20+E | 934 | W0 DATA | TCCl0.12_V_1 te=te:20 scalarw(3) @_SINT/CC/MAPR10NoCE1_ARA0 te=te:20 write(0, 0) |
//| 35   | 934 | W1 DATA |                                                                                  |
//| 20   | 935 | R0 DATA |                                                                                  |
//| 20+E | 935 | W0 DATA | TCCl0.12_V_1 te=te:20 scalarw(3) @_SINT/CC/MAPR10NoCE0_ARA0 te=te:20 write(0, 0) |
//| 36   | 935 | W1 DATA |                                                                                  |
//| 20   | 936 | R0 DATA |                                                                                  |
//| 20+E | 936 | W0 DATA | TCCl0.12_V_1 te=te:20 scalarw(4) TCCl0.12_V_0 te=te:20 scalarw(1+TCCl0.12_V_0)   |
//*------+-----+---------+----------------------------------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X21:"xpc10:21" 949 :  major_start_pcl=37   edge_private_start/end=-1/-1 exec=37 (dend=0)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X21:"xpc10:21" 948 :  major_start_pcl=37   edge_private_start/end=49/49 exec=37 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X21:"xpc10:21" 947 :  major_start_pcl=37   edge_private_start/end=48/48 exec=37 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X21:"xpc10:21" 946 :  major_start_pcl=37   edge_private_start/end=47/47 exec=37 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X21:"xpc10:21" 945 :  major_start_pcl=37   edge_private_start/end=46/46 exec=37 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X21:"xpc10:21" 944 :  major_start_pcl=37   edge_private_start/end=45/45 exec=37 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X21:"xpc10:21" 943 :  major_start_pcl=37   edge_private_start/end=44/44 exec=37 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X21:"xpc10:21" 942 :  major_start_pcl=37   edge_private_start/end=43/43 exec=37 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X21:"xpc10:21" 941 :  major_start_pcl=37   edge_private_start/end=42/42 exec=37 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X21:"xpc10:21" 940 :  major_start_pcl=37   edge_private_start/end=41/41 exec=37 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X21:"xpc10:21" 939 :  major_start_pcl=37   edge_private_start/end=40/40 exec=37 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X21:"xpc10:21" 938 :  major_start_pcl=37   edge_private_start/end=39/39 exec=37 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X21:"xpc10:21" 937 :  major_start_pcl=37   edge_private_start/end=38/38 exec=37 (dend=1)
//Simple greedy schedule for res2: Thread=xpc10 state=X21:"xpc10:21"
//res2: Thread=xpc10 state=X21:"xpc10:21"
//*------+-----+---------+----------------------------------------------------------------------------------*
//| pc   | eno | Phaser  | Work                                                                             |
//*------+-----+---------+----------------------------------------------------------------------------------*
//| 37   | -   | R0 CTRL |                                                                                  |
//| 37   | 937 | R0 DATA |                                                                                  |
//| 37+E | 937 | W0 DATA | TCCl0.12_V_1 te=te:37 scalarw(2) @_SINT/CC/MAPR10NoCE3_ARA0 te=te:37 write(0, 0) |
//| 38   | 937 | W1 DATA |                                                                                  |
//| 37   | 938 | R0 DATA |                                                                                  |
//| 37+E | 938 | W0 DATA | TCCl0.12_V_1 te=te:37 scalarw(2) @_SINT/CC/MAPR10NoCE2_ARA0 te=te:37 write(0, 0) |
//| 39   | 938 | W1 DATA |                                                                                  |
//| 37   | 939 | R0 DATA |                                                                                  |
//| 37+E | 939 | W0 DATA | TCCl0.12_V_1 te=te:37 scalarw(2) @_SINT/CC/MAPR10NoCE1_ARA0 te=te:37 write(0, 0) |
//| 40   | 939 | W1 DATA |                                                                                  |
//| 37   | 940 | R0 DATA |                                                                                  |
//| 37+E | 940 | W0 DATA | TCCl0.12_V_1 te=te:37 scalarw(2) @_SINT/CC/MAPR10NoCE0_ARA0 te=te:37 write(0, 0) |
//| 41   | 940 | W1 DATA |                                                                                  |
//| 37   | 941 | R0 DATA |                                                                                  |
//| 37+E | 941 | W0 DATA | TCCl0.12_V_1 te=te:37 scalarw(2) @_SINT/CC/MAPR10NoCE3_ARA0 te=te:37 write(0, 0) |
//| 42   | 941 | W1 DATA |                                                                                  |
//| 37   | 942 | R0 DATA |                                                                                  |
//| 37+E | 942 | W0 DATA | TCCl0.12_V_1 te=te:37 scalarw(2) @_SINT/CC/MAPR10NoCE2_ARA0 te=te:37 write(0, 0) |
//| 43   | 942 | W1 DATA |                                                                                  |
//| 37   | 943 | R0 DATA |                                                                                  |
//| 37+E | 943 | W0 DATA | TCCl0.12_V_1 te=te:37 scalarw(2) @_SINT/CC/MAPR10NoCE1_ARA0 te=te:37 write(0, 0) |
//| 44   | 943 | W1 DATA |                                                                                  |
//| 37   | 944 | R0 DATA |                                                                                  |
//| 37+E | 944 | W0 DATA | TCCl0.12_V_1 te=te:37 scalarw(2) @_SINT/CC/MAPR10NoCE0_ARA0 te=te:37 write(0, 0) |
//| 45   | 944 | W1 DATA |                                                                                  |
//| 37   | 945 | R0 DATA |                                                                                  |
//| 37+E | 945 | W0 DATA | TCCl0.12_V_1 te=te:37 scalarw(3) @_SINT/CC/MAPR10NoCE3_ARA0 te=te:37 write(0, 0) |
//| 46   | 945 | W1 DATA |                                                                                  |
//| 37   | 946 | R0 DATA |                                                                                  |
//| 37+E | 946 | W0 DATA | TCCl0.12_V_1 te=te:37 scalarw(3) @_SINT/CC/MAPR10NoCE2_ARA0 te=te:37 write(0, 0) |
//| 47   | 946 | W1 DATA |                                                                                  |
//| 37   | 947 | R0 DATA |                                                                                  |
//| 37+E | 947 | W0 DATA | TCCl0.12_V_1 te=te:37 scalarw(3) @_SINT/CC/MAPR10NoCE1_ARA0 te=te:37 write(0, 0) |
//| 48   | 947 | W1 DATA |                                                                                  |
//| 37   | 948 | R0 DATA |                                                                                  |
//| 37+E | 948 | W0 DATA | TCCl0.12_V_1 te=te:37 scalarw(3) @_SINT/CC/MAPR10NoCE0_ARA0 te=te:37 write(0, 0) |
//| 49   | 948 | W1 DATA |                                                                                  |
//| 37   | 949 | R0 DATA |                                                                                  |
//| 37+E | 949 | W0 DATA | TCCl0.12_V_1 te=te:37 scalarw(4) TCCl0.12_V_0 te=te:37 scalarw(1+TCCl0.12_V_0)   |
//*------+-----+---------+----------------------------------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X22:"xpc10:22" 958 :  major_start_pcl=50   edge_private_start/end=-1/-1 exec=50 (dend=0)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X22:"xpc10:22" 957 :  major_start_pcl=50   edge_private_start/end=58/58 exec=50 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X22:"xpc10:22" 956 :  major_start_pcl=50   edge_private_start/end=57/57 exec=50 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X22:"xpc10:22" 955 :  major_start_pcl=50   edge_private_start/end=56/56 exec=50 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X22:"xpc10:22" 954 :  major_start_pcl=50   edge_private_start/end=55/55 exec=50 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X22:"xpc10:22" 953 :  major_start_pcl=50   edge_private_start/end=54/54 exec=50 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X22:"xpc10:22" 952 :  major_start_pcl=50   edge_private_start/end=53/53 exec=50 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X22:"xpc10:22" 951 :  major_start_pcl=50   edge_private_start/end=52/52 exec=50 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X22:"xpc10:22" 950 :  major_start_pcl=50   edge_private_start/end=51/51 exec=50 (dend=1)
//Simple greedy schedule for res2: Thread=xpc10 state=X22:"xpc10:22"
//res2: Thread=xpc10 state=X22:"xpc10:22"
//*------+-----+---------+----------------------------------------------------------------------------------*
//| pc   | eno | Phaser  | Work                                                                             |
//*------+-----+---------+----------------------------------------------------------------------------------*
//| 50   | -   | R0 CTRL |                                                                                  |
//| 50   | 950 | R0 DATA |                                                                                  |
//| 50+E | 950 | W0 DATA | TCCl0.12_V_1 te=te:50 scalarw(3) @_SINT/CC/MAPR10NoCE3_ARA0 te=te:50 write(0, 0) |
//| 51   | 950 | W1 DATA |                                                                                  |
//| 50   | 951 | R0 DATA |                                                                                  |
//| 50+E | 951 | W0 DATA | TCCl0.12_V_1 te=te:50 scalarw(3) @_SINT/CC/MAPR10NoCE2_ARA0 te=te:50 write(0, 0) |
//| 52   | 951 | W1 DATA |                                                                                  |
//| 50   | 952 | R0 DATA |                                                                                  |
//| 50+E | 952 | W0 DATA | TCCl0.12_V_1 te=te:50 scalarw(3) @_SINT/CC/MAPR10NoCE1_ARA0 te=te:50 write(0, 0) |
//| 53   | 952 | W1 DATA |                                                                                  |
//| 50   | 953 | R0 DATA |                                                                                  |
//| 50+E | 953 | W0 DATA | TCCl0.12_V_1 te=te:50 scalarw(3) @_SINT/CC/MAPR10NoCE0_ARA0 te=te:50 write(0, 0) |
//| 54   | 953 | W1 DATA |                                                                                  |
//| 50   | 954 | R0 DATA |                                                                                  |
//| 50+E | 954 | W0 DATA | TCCl0.12_V_1 te=te:50 scalarw(3) @_SINT/CC/MAPR10NoCE3_ARA0 te=te:50 write(0, 0) |
//| 55   | 954 | W1 DATA |                                                                                  |
//| 50   | 955 | R0 DATA |                                                                                  |
//| 50+E | 955 | W0 DATA | TCCl0.12_V_1 te=te:50 scalarw(3) @_SINT/CC/MAPR10NoCE2_ARA0 te=te:50 write(0, 0) |
//| 56   | 955 | W1 DATA |                                                                                  |
//| 50   | 956 | R0 DATA |                                                                                  |
//| 50+E | 956 | W0 DATA | TCCl0.12_V_1 te=te:50 scalarw(3) @_SINT/CC/MAPR10NoCE1_ARA0 te=te:50 write(0, 0) |
//| 57   | 956 | W1 DATA |                                                                                  |
//| 50   | 957 | R0 DATA |                                                                                  |
//| 50+E | 957 | W0 DATA | TCCl0.12_V_1 te=te:50 scalarw(3) @_SINT/CC/MAPR10NoCE0_ARA0 te=te:50 write(0, 0) |
//| 58   | 957 | W1 DATA |                                                                                  |
//| 50   | 958 | R0 DATA |                                                                                  |
//| 50+E | 958 | W0 DATA | TCCl0.12_V_1 te=te:50 scalarw(4) TCCl0.12_V_0 te=te:50 scalarw(1+TCCl0.12_V_0)   |
//*------+-----+---------+----------------------------------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X23:"xpc10:23" 963 :  major_start_pcl=59   edge_private_start/end=-1/-1 exec=59 (dend=0)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X23:"xpc10:23" 962 :  major_start_pcl=59   edge_private_start/end=63/63 exec=59 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X23:"xpc10:23" 961 :  major_start_pcl=59   edge_private_start/end=62/62 exec=59 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X23:"xpc10:23" 960 :  major_start_pcl=59   edge_private_start/end=61/61 exec=59 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X23:"xpc10:23" 959 :  major_start_pcl=59   edge_private_start/end=60/60 exec=59 (dend=1)
//Simple greedy schedule for res2: Thread=xpc10 state=X23:"xpc10:23"
//res2: Thread=xpc10 state=X23:"xpc10:23"
//*------+-----+---------+----------------------------------------------------------------------------------*
//| pc   | eno | Phaser  | Work                                                                             |
//*------+-----+---------+----------------------------------------------------------------------------------*
//| 59   | -   | R0 CTRL |                                                                                  |
//| 59   | 959 | R0 DATA |                                                                                  |
//| 59+E | 959 | W0 DATA | TCCl0.12_V_1 te=te:59 scalarw(4) @_SINT/CC/MAPR10NoCE3_ARA0 te=te:59 write(0, 0) |
//| 60   | 959 | W1 DATA |                                                                                  |
//| 59   | 960 | R0 DATA |                                                                                  |
//| 59+E | 960 | W0 DATA | TCCl0.12_V_1 te=te:59 scalarw(4) @_SINT/CC/MAPR10NoCE2_ARA0 te=te:59 write(0, 0) |
//| 61   | 960 | W1 DATA |                                                                                  |
//| 59   | 961 | R0 DATA |                                                                                  |
//| 59+E | 961 | W0 DATA | TCCl0.12_V_1 te=te:59 scalarw(4) @_SINT/CC/MAPR10NoCE1_ARA0 te=te:59 write(0, 0) |
//| 62   | 961 | W1 DATA |                                                                                  |
//| 59   | 962 | R0 DATA |                                                                                  |
//| 59+E | 962 | W0 DATA | TCCl0.12_V_1 te=te:59 scalarw(4) @_SINT/CC/MAPR10NoCE0_ARA0 te=te:59 write(0, 0) |
//| 63   | 962 | W1 DATA |                                                                                  |
//| 59   | 963 | R0 DATA |                                                                                  |
//| 59+E | 963 | W0 DATA | TCCl0.12_V_1 te=te:59 scalarw(4) TCCl0.12_V_0 te=te:59 scalarw(1+TCCl0.12_V_0)   |
//*------+-----+---------+----------------------------------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X24:"xpc10:24" 964 :  major_start_pcl=64   edge_private_start/end=-1/-1 exec=64 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X24:"xpc10:24"
//res2: Thread=xpc10 state=X24:"xpc10:24"
//*------+-----+---------+-----------------------------------------------*
//| pc   | eno | Phaser  | Work                                          |
//*------+-----+---------+-----------------------------------------------*
//| 64   | -   | R0 CTRL |                                               |
//| 64   | 964 | R0 DATA |                                               |
//| 64+E | 964 | W0 DATA | TCCl0.12_V_0 te=te:64 scalarw(1+TCCl0.12_V_0) |
//*------+-----+---------+-----------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X25:"xpc10:25" 982 :  major_start_pcl=65   edge_private_start/end=81/81 exec=65 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X25:"xpc10:25" 981 :  major_start_pcl=65   edge_private_start/end=80/80 exec=65 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X25:"xpc10:25" 980 :  major_start_pcl=65   edge_private_start/end=79/79 exec=65 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X25:"xpc10:25" 979 :  major_start_pcl=65   edge_private_start/end=78/78 exec=65 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X25:"xpc10:25" 978 :  major_start_pcl=65   edge_private_start/end=77/77 exec=65 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X25:"xpc10:25" 977 :  major_start_pcl=65   edge_private_start/end=76/76 exec=65 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X25:"xpc10:25" 976 :  major_start_pcl=65   edge_private_start/end=75/75 exec=65 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X25:"xpc10:25" 975 :  major_start_pcl=65   edge_private_start/end=74/74 exec=65 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X25:"xpc10:25" 974 :  major_start_pcl=65   edge_private_start/end=73/73 exec=65 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X25:"xpc10:25" 973 :  major_start_pcl=65   edge_private_start/end=72/72 exec=65 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X25:"xpc10:25" 972 :  major_start_pcl=65   edge_private_start/end=71/71 exec=65 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X25:"xpc10:25" 971 :  major_start_pcl=65   edge_private_start/end=70/70 exec=65 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X25:"xpc10:25" 970 :  major_start_pcl=65   edge_private_start/end=69/69 exec=65 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X25:"xpc10:25" 969 :  major_start_pcl=65   edge_private_start/end=68/68 exec=65 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X25:"xpc10:25" 968 :  major_start_pcl=65   edge_private_start/end=67/67 exec=65 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X25:"xpc10:25" 967 :  major_start_pcl=65   edge_private_start/end=66/66 exec=65 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X25:"xpc10:25" 966 :  major_start_pcl=65   edge_private_start/end=-1/-1 exec=65 (dend=0)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X25:"xpc10:25" 965 :  major_start_pcl=65   edge_private_start/end=-1/-1 exec=65 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X25:"xpc10:25"
//res2: Thread=xpc10 state=X25:"xpc10:25"
//*------+-----+---------+---------------------------------------------------------------------------------------------*
//| pc   | eno | Phaser  | Work                                                                                        |
//*------+-----+---------+---------------------------------------------------------------------------------------------*
//| 65   | -   | R0 CTRL |                                                                                             |
//| 65   | 965 | R0 DATA |                                                                                             |
//| 65+E | 965 | W0 DATA | TCCl0.12_V_1 te=te:65 scalarw(4) TCCl0.12_V_0 te=te:65 scalarw(1+TCCl0.12_V_0)              |
//| 65   | 966 | R0 DATA |                                                                                             |
//| 65+E | 966 | W0 DATA |  W/P:Cache Cleared  PLI:Cuckoo cache cleared                                                |
//| 65   | 967 | R0 DATA |                                                                                             |
//| 65+E | 967 | W0 DATA | TCCl0.12_V_1 te=te:65 scalarw(0) @_SINT/CC/MAPR10NoCE3_ARA0 te=te:65 write(TCCl0.12_V_0, 0) |
//| 66   | 967 | W1 DATA |                                                                                             |
//| 65   | 968 | R0 DATA |                                                                                             |
//| 65+E | 968 | W0 DATA | TCCl0.12_V_1 te=te:65 scalarw(0) @_SINT/CC/MAPR10NoCE2_ARA0 te=te:65 write(TCCl0.12_V_0, 0) |
//| 67   | 968 | W1 DATA |                                                                                             |
//| 65   | 969 | R0 DATA |                                                                                             |
//| 65+E | 969 | W0 DATA | TCCl0.12_V_1 te=te:65 scalarw(0) @_SINT/CC/MAPR10NoCE1_ARA0 te=te:65 write(TCCl0.12_V_0, 0) |
//| 68   | 969 | W1 DATA |                                                                                             |
//| 65   | 970 | R0 DATA |                                                                                             |
//| 65+E | 970 | W0 DATA | TCCl0.12_V_1 te=te:65 scalarw(0) @_SINT/CC/MAPR10NoCE0_ARA0 te=te:65 write(TCCl0.12_V_0, 0) |
//| 69   | 970 | W1 DATA |                                                                                             |
//| 65   | 971 | R0 DATA |                                                                                             |
//| 65+E | 971 | W0 DATA | TCCl0.12_V_1 te=te:65 scalarw(1) @_SINT/CC/MAPR10NoCE3_ARA0 te=te:65 write(TCCl0.12_V_0, 0) |
//| 70   | 971 | W1 DATA |                                                                                             |
//| 65   | 972 | R0 DATA |                                                                                             |
//| 65+E | 972 | W0 DATA | TCCl0.12_V_1 te=te:65 scalarw(1) @_SINT/CC/MAPR10NoCE2_ARA0 te=te:65 write(TCCl0.12_V_0, 0) |
//| 71   | 972 | W1 DATA |                                                                                             |
//| 65   | 973 | R0 DATA |                                                                                             |
//| 65+E | 973 | W0 DATA | TCCl0.12_V_1 te=te:65 scalarw(1) @_SINT/CC/MAPR10NoCE1_ARA0 te=te:65 write(TCCl0.12_V_0, 0) |
//| 72   | 973 | W1 DATA |                                                                                             |
//| 65   | 974 | R0 DATA |                                                                                             |
//| 65+E | 974 | W0 DATA | TCCl0.12_V_1 te=te:65 scalarw(1) @_SINT/CC/MAPR10NoCE0_ARA0 te=te:65 write(TCCl0.12_V_0, 0) |
//| 73   | 974 | W1 DATA |                                                                                             |
//| 65   | 975 | R0 DATA |                                                                                             |
//| 65+E | 975 | W0 DATA | TCCl0.12_V_1 te=te:65 scalarw(2) @_SINT/CC/MAPR10NoCE3_ARA0 te=te:65 write(TCCl0.12_V_0, 0) |
//| 74   | 975 | W1 DATA |                                                                                             |
//| 65   | 976 | R0 DATA |                                                                                             |
//| 65+E | 976 | W0 DATA | TCCl0.12_V_1 te=te:65 scalarw(2) @_SINT/CC/MAPR10NoCE2_ARA0 te=te:65 write(TCCl0.12_V_0, 0) |
//| 75   | 976 | W1 DATA |                                                                                             |
//| 65   | 977 | R0 DATA |                                                                                             |
//| 65+E | 977 | W0 DATA | TCCl0.12_V_1 te=te:65 scalarw(2) @_SINT/CC/MAPR10NoCE1_ARA0 te=te:65 write(TCCl0.12_V_0, 0) |
//| 76   | 977 | W1 DATA |                                                                                             |
//| 65   | 978 | R0 DATA |                                                                                             |
//| 65+E | 978 | W0 DATA | TCCl0.12_V_1 te=te:65 scalarw(2) @_SINT/CC/MAPR10NoCE0_ARA0 te=te:65 write(TCCl0.12_V_0, 0) |
//| 77   | 978 | W1 DATA |                                                                                             |
//| 65   | 979 | R0 DATA |                                                                                             |
//| 65+E | 979 | W0 DATA | TCCl0.12_V_1 te=te:65 scalarw(3) @_SINT/CC/MAPR10NoCE3_ARA0 te=te:65 write(TCCl0.12_V_0, 0) |
//| 78   | 979 | W1 DATA |                                                                                             |
//| 65   | 980 | R0 DATA |                                                                                             |
//| 65+E | 980 | W0 DATA | TCCl0.12_V_1 te=te:65 scalarw(3) @_SINT/CC/MAPR10NoCE2_ARA0 te=te:65 write(TCCl0.12_V_0, 0) |
//| 79   | 980 | W1 DATA |                                                                                             |
//| 65   | 981 | R0 DATA |                                                                                             |
//| 65+E | 981 | W0 DATA | TCCl0.12_V_1 te=te:65 scalarw(3) @_SINT/CC/MAPR10NoCE1_ARA0 te=te:65 write(TCCl0.12_V_0, 0) |
//| 80   | 981 | W1 DATA |                                                                                             |
//| 65   | 982 | R0 DATA |                                                                                             |
//| 65+E | 982 | W0 DATA | TCCl0.12_V_1 te=te:65 scalarw(3) @_SINT/CC/MAPR10NoCE0_ARA0 te=te:65 write(TCCl0.12_V_0, 0) |
//| 81   | 982 | W1 DATA |                                                                                             |
//*------+-----+---------+---------------------------------------------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X26:"xpc10:26" 983 :  major_start_pcl=82   edge_private_start/end=-1/-1 exec=82 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X26:"xpc10:26"
//res2: Thread=xpc10 state=X26:"xpc10:26"
//*------+-----+---------+---------------------------------------------------------------------------------------------------------------------*
//| pc   | eno | Phaser  | Work                                                                                                                |
//*------+-----+---------+---------------------------------------------------------------------------------------------------------------------*
//| 82   | -   | R0 CTRL |                                                                                                                     |
//| 82   | 983 | R0 DATA |                                                                                                                     |
//| 82+E | 983 | W0 DATA | @64_US/CC/SCALbx28_dk te=te:82 scalarw(U64'9999999900000000I) @_SINT/CC/SCALbx28_seed te=te:82 scalarw(S32'123456I) |
//*------+-----+---------+---------------------------------------------------------------------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X27:"xpc10:27" 984 :  major_start_pcl=83   edge_private_start/end=-1/-1 exec=83 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X27:"xpc10:27"
//res2: Thread=xpc10 state=X27:"xpc10:27"
//*------+-----+---------+-------------------------------------------------------*
//| pc   | eno | Phaser  | Work                                                  |
//*------+-----+---------+-------------------------------------------------------*
//| 83   | -   | R0 CTRL |                                                       |
//| 83   | 984 | R0 DATA |                                                       |
//| 83+E | 984 | W0 DATA | @_SINT/CC/SCALbx28_seed te=te:83 scalarw(S32'123456I) |
//*------+-----+---------+-------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X28:"xpc10:28" 985 :  major_start_pcl=84   edge_private_start/end=-1/-1 exec=84 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X28:"xpc10:28"
//res2: Thread=xpc10 state=X28:"xpc10:28"
//*------+-----+---------+-------------------------------------------------------------------------------------------------*
//| pc   | eno | Phaser  | Work                                                                                            |
//*------+-----+---------+-------------------------------------------------------------------------------------------------*
//| 84   | -   | R0 CTRL |                                                                                                 |
//| 84   | 985 | R0 DATA |                                                                                                 |
//| 84+E | 985 | W0 DATA | @64_US/CC/SCALbx28_dk te=te:84 scalarw(U64'9999999900000000I) TTMT4Main_V_2 te=te:84 scalarw(0) |
//*------+-----+---------+-------------------------------------------------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X29:"xpc10:29" 986 :  major_start_pcl=85   edge_private_start/end=-1/-1 exec=85 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X29:"xpc10:29"
//res2: Thread=xpc10 state=X29:"xpc10:29"
//*------+-----+---------+---------------------------------------------------------------------*
//| pc   | eno | Phaser  | Work                                                                |
//*------+-----+---------+---------------------------------------------------------------------*
//| 85   | -   | R0 CTRL |                                                                     |
//| 85   | 986 | R0 DATA |                                                                     |
//| 85+E | 986 | W0 DATA | TTMT4Main_V_4 te=te:85 scalarw(0) TTMT4Main_V_3 te=te:85 scalarw(0) |
//*------+-----+---------+---------------------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X30:"xpc10:30" 988 :  major_start_pcl=86   edge_private_start/end=-1/-1 exec=86 (dend=0)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X30:"xpc10:30" 987 :  major_start_pcl=86   edge_private_start/end=-1/-1 exec=86 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X30:"xpc10:30"
//res2: Thread=xpc10 state=X30:"xpc10:30"
//*------+-----+---------+------------------------------------------------*
//| pc   | eno | Phaser  | Work                                           |
//*------+-----+---------+------------------------------------------------*
//| 86   | -   | R0 CTRL |                                                |
//| 86   | 987 | R0 DATA |                                                |
//| 86+E | 987 | W0 DATA |  W/P:Data Entered  PLI:Cuckoo cache inserte... |
//| 86   | 988 | R0 DATA |                                                |
//| 86+E | 988 | W0 DATA | @_SINT/CC/SCALbx28_seed te=te:86 scalarw(E1)   |
//*------+-----+---------+------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X31:"xpc10:31" 989 :  major_start_pcl=87   edge_private_start/end=-1/-1 exec=87 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X31:"xpc10:31"
//res2: Thread=xpc10 state=X31:"xpc10:31"
//*------+-----+---------+---------------------------------------------------------------------------------------------------------------------*
//| pc   | eno | Phaser  | Work                                                                                                                |
//*------+-----+---------+---------------------------------------------------------------------------------------------------------------------*
//| 87   | -   | R0 CTRL |                                                                                                                     |
//| 87   | 989 | R0 DATA |                                                                                                                     |
//| 87+E | 989 | W0 DATA | @64_US/CC/SCALbx28_dk te=te:87 scalarw(U64'9999999900000000I) @_SINT/CC/SCALbx28_seed te=te:87 scalarw(S32'123456I) |
//*------+-----+---------+---------------------------------------------------------------------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X32:"xpc10:32" 990 :  major_start_pcl=88   edge_private_start/end=-1/-1 exec=88 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X32:"xpc10:32"
//res2: Thread=xpc10 state=X32:"xpc10:32"
//*------+-----+---------+---------------------------------------------------------------------*
//| pc   | eno | Phaser  | Work                                                                |
//*------+-----+---------+---------------------------------------------------------------------*
//| 88   | -   | R0 CTRL |                                                                     |
//| 88   | 990 | R0 DATA |                                                                     |
//| 88+E | 990 | W0 DATA | TTMT4Main_V_9 te=te:88 scalarw(0) TTMT4Main_V_8 te=te:88 scalarw(0) |
//*------+-----+---------+---------------------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X33:"xpc10:33" 991 :  major_start_pcl=89   edge_private_start/end=-1/-1 exec=89 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X33:"xpc10:33"
//res2: Thread=xpc10 state=X33:"xpc10:33"
//*------+-----+---------+---------------------------------------------------------------------------------*
//| pc   | eno | Phaser  | Work                                                                            |
//*------+-----+---------+---------------------------------------------------------------------------------*
//| 89   | -   | R0 CTRL |                                                                                 |
//| 89   | 991 | R0 DATA |                                                                                 |
//| 89+E | 991 | W0 DATA | @_SINT/CC/SCALbx28_seed te=te:89 scalarw(E1) TTMT4Main_V_10 te=te:89 scalarw(0) |
//*------+-----+---------+---------------------------------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X34:"xpc10:34" 992 :  major_start_pcl=90   edge_private_start/end=-1/-1 exec=90 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X34:"xpc10:34"
//res2: Thread=xpc10 state=X34:"xpc10:34"
//*------+-----+---------+-------------------------------------*
//| pc   | eno | Phaser  | Work                                |
//*------+-----+---------+-------------------------------------*
//| 90   | -   | R0 CTRL |                                     |
//| 90   | 992 | R0 DATA |                                     |
//| 90+E | 992 | W0 DATA | TTMT4Main_V_11 te=te:90 scalarw(E2) |
//*------+-----+---------+-------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X35:"xpc10:35" 993 :  major_start_pcl=91   edge_private_start/end=-1/-1 exec=91 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X35:"xpc10:35"
//res2: Thread=xpc10 state=X35:"xpc10:35"
//*------+-----+---------+----------------------------------------------------------------------*
//| pc   | eno | Phaser  | Work                                                                 |
//*------+-----+---------+----------------------------------------------------------------------*
//| 91   | -   | R0 CTRL |                                                                      |
//| 91   | 993 | R0 DATA |                                                                      |
//| 91+E | 993 | W0 DATA | TDGe6.4_V_0 te=te:91 scalarw(E3) fastspilldup30 te=te:91 scalarw(E3) |
//*------+-----+---------+----------------------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X36:"xpc10:36" 994 :  major_start_pcl=92   edge_private_start/end=-1/-1 exec=92 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X36:"xpc10:36"
//res2: Thread=xpc10 state=X36:"xpc10:36"
//*------+-----+---------+---------------------------------------------------------------*
//| pc   | eno | Phaser  | Work                                                          |
//*------+-----+---------+---------------------------------------------------------------*
//| 92   | -   | R0 CTRL |                                                               |
//| 92   | 994 | R0 DATA |                                                               |
//| 92+E | 994 | W0 DATA | @64_US/CC/SCALbx28_dk te=te:92 scalarw(S64'1I+fastspilldup30) |
//*------+-----+---------+---------------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X37:"xpc10:37" 995 :  major_start_pcl=93   edge_private_start/end=-1/-1 exec=93 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X37:"xpc10:37"
//res2: Thread=xpc10 state=X37:"xpc10:37"
//*------+-----+---------+----------------------------------------------------*
//| pc   | eno | Phaser  | Work                                               |
//*------+-----+---------+----------------------------------------------------*
//| 93   | -   | R0 CTRL |                                                    |
//| 93   | 995 | R0 DATA |                                                    |
//| 93+E | 995 | W0 DATA | TTMT4Main_V_12 te=te:93 scalarw(C64u(TDGe6.4_V_0)) |
//*------+-----+---------+----------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X38:"xpc10:38" 996 :  major_start_pcl=94   edge_private_start/end=-1/-1 exec=94 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X38:"xpc10:38"
//res2: Thread=xpc10 state=X38:"xpc10:38"
//*------+-----+---------+-------------------------------------------------------*
//| pc   | eno | Phaser  | Work                                                  |
//*------+-----+---------+-------------------------------------------------------*
//| 94   | -   | R0 CTRL |                                                       |
//| 94   | 996 | R0 DATA |                                                       |
//| 94+E | 996 | W0 DATA | @_SINT/CC/SCALbx24_stats_lookups te=te:94 scalarw(E4) |
//*------+-----+---------+-------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X39:"xpc10:39" 998 :  major_start_pcl=95   edge_private_start/end=-1/-1 exec=95 (dend=0)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X39:"xpc10:39" 997 :  major_start_pcl=95   edge_private_start/end=-1/-1 exec=95 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X39:"xpc10:39"
//res2: Thread=xpc10 state=X39:"xpc10:39"
//*------+-----+---------+------------------------------------------------------------------------------*
//| pc   | eno | Phaser  | Work                                                                         |
//*------+-----+---------+------------------------------------------------------------------------------*
//| 95   | -   | R0 CTRL |                                                                              |
//| 95   | 997 | R0 DATA |                                                                              |
//| 95+E | 997 | W0 DATA | TCl6._SPILL_256 te=te:95 scalarw(-4) TTMT4Main_V_13 te=te:95 scalarw(U64'0I) |
//| 95   | 998 | R0 DATA |                                                                              |
//| 95+E | 998 | W0 DATA | TTMT4Main_V_13 te=te:95 scalarw(U64'0I) TClo6.9_V_1 te=te:95 scalarw(0)      |
//*------+-----+---------+------------------------------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X40:"xpc10:40" 1001 :  major_start_pcl=96   edge_private_start/end=-1/-1 exec=96 (dend=0)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X40:"xpc10:40" 1000 :  major_start_pcl=96   edge_private_start/end=-1/-1 exec=96 (dend=0)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X40:"xpc10:40" 999 :  major_start_pcl=96   edge_private_start/end=-1/-1 exec=96 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X40:"xpc10:40"
//res2: Thread=xpc10 state=X40:"xpc10:40"
//*------+------+---------+-----------------------------------------------------------------------------------------------------*
//| pc   | eno  | Phaser  | Work                                                                                                |
//*------+------+---------+-----------------------------------------------------------------------------------------------------*
//| 96   | -    | R0 CTRL |                                                                                                     |
//| 96   | 999  | R0 DATA |                                                                                                     |
//| 96+E | 999  | W0 DATA | TTMT4Main_V_9 te=te:96 scalarw(1+TTMT4Main_V_9) TTMT4Main_V_14 te=te:96 scalarw(C(TCl6._SPILL_256)) |
//| 96   | 1000 | R0 DATA |                                                                                                     |
//| 96+E | 1000 | W0 DATA | TTMT4Main_V_8 te=te:96 scalarw(1+TTMT4Main_V_8) TTMT4Main_V_14 te=te:96 scalarw(C(TCl6._SPILL_256)) |
//| 96   | 1001 | R0 DATA |                                                                                                     |
//| 96+E | 1001 | W0 DATA | TTMT4Main_V_8 te=te:96 scalarw(1+TTMT4Main_V_8) TTMT4Main_V_14 te=te:96 scalarw(C(TCl6._SPILL_256)) |
//*------+------+---------+-----------------------------------------------------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X41:"xpc10:41" 1002 :  major_start_pcl=97   edge_private_start/end=-1/-1 exec=97 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X41:"xpc10:41"
//res2: Thread=xpc10 state=X41:"xpc10:41"
//*------+------+---------+-------------------------------------------------*
//| pc   | eno  | Phaser  | Work                                            |
//*------+------+---------+-------------------------------------------------*
//| 97   | -    | R0 CTRL |                                                 |
//| 97   | 1002 | R0 DATA |                                                 |
//| 97+E | 1002 | W0 DATA | TTMT4Main_V_8 te=te:97 scalarw(1+TTMT4Main_V_8) |
//*------+------+---------+-------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X42:"xpc10:42" 1003 :  major_start_pcl=98   edge_private_start/end=-1/-1 exec=98 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X42:"xpc10:42"
//res2: Thread=xpc10 state=X42:"xpc10:42"
//*------+------+---------+---------------------------------------------------*
//| pc   | eno  | Phaser  | Work                                              |
//*------+------+---------+---------------------------------------------------*
//| 98   | -    | R0 CTRL |                                                   |
//| 98   | 1003 | R0 DATA |                                                   |
//| 98+E | 1003 | W0 DATA | TTMT4Main_V_10 te=te:98 scalarw(1+TTMT4Main_V_10) |
//*------+------+---------+---------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X43:"xpc10:43" 1005 :  major_start_pcl=99   edge_private_start/end=-1/-1 exec=99 (dend=0)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X43:"xpc10:43" 1004 :  major_start_pcl=99   edge_private_start/end=-1/-1 exec=99 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X43:"xpc10:43"
//res2: Thread=xpc10 state=X43:"xpc10:43"
//*------+------+---------+-------------------------------------------------*
//| pc   | eno  | Phaser  | Work                                            |
//*------+------+---------+-------------------------------------------------*
//| 99   | -    | R0 CTRL |                                                 |
//| 99   | 1004 | R0 DATA |                                                 |
//| 99+E | 1004 | W0 DATA |  W/P:Readback Done  PLI:Cuckoo cache inserte... |
//| 99   | 1005 | R0 DATA |                                                 |
//| 99+E | 1005 | W0 DATA | @_SINT/CC/SCALbx28_seed te=te:99 scalarw(E1)    |
//*------+------+---------+-------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X44:"xpc10:44" 1006 :  major_start_pcl=100   edge_private_start/end=-1/-1 exec=100 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X44:"xpc10:44"
//res2: Thread=xpc10 state=X44:"xpc10:44"
//*-------+------+---------+-----------------------------------------------------------*
//| pc    | eno  | Phaser  | Work                                                      |
//*-------+------+---------+-----------------------------------------------------------*
//| 100   | -    | R0 CTRL |                                                           |
//| 100   | 1006 | R0 DATA |                                                           |
//| 100+E | 1006 | W0 DATA |  PLI:cuckoo cache: insert...  PLI:cuckoo cache: this=%... |
//*-------+------+---------+-----------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X45:"xpc10:45" 1007 :  major_start_pcl=101   edge_private_start/end=-1/-1 exec=101 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X45:"xpc10:45"
//res2: Thread=xpc10 state=X45:"xpc10:45"
//*-------+------+---------+-----------------------------------------------------------*
//| pc    | eno  | Phaser  | Work                                                      |
//*-------+------+---------+-----------------------------------------------------------*
//| 101   | -    | R0 CTRL |                                                           |
//| 101   | 1007 | R0 DATA |                                                           |
//| 101+E | 1007 | W0 DATA |  PLI:Cuckoo cache demo fi...  PLI:cuckoo cache: lookup... |
//*-------+------+---------+-----------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X46:"xpc10:46" 1008 :  major_start_pcl=102   edge_private_start/end=-1/-1 exec=102 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X46:"xpc10:46"
//res2: Thread=xpc10 state=X46:"xpc10:46"
//*-------+------+---------+-----------------------------------------------------*
//| pc    | eno  | Phaser  | Work                                                |
//*-------+------+---------+-----------------------------------------------------*
//| 102   | -    | R0 CTRL |                                                     |
//| 102   | 1008 | R0 DATA |                                                     |
//| 102+E | 1008 | W0 DATA | done te=te:102 scalarw(U1'1I)  PLI:GSAI:hpr_sysexit |
//*-------+------+---------+-----------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X47:"xpc10:47" 1009 :  major_start_pcl=103   edge_private_start/end=-1/-1 exec=103 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X47:"xpc10:47"
//res2: Thread=xpc10 state=X47:"xpc10:47"
//*-------+------+---------+----------------------------------*
//| pc    | eno  | Phaser  | Work                             |
//*-------+------+---------+----------------------------------*
//| 103   | -    | R0 CTRL |                                  |
//| 103   | 1009 | R0 DATA |                                  |
//| 103+E | 1009 | W0 DATA | TClo6.9_V_0 te=te:103 scalarw(0) |
//*-------+------+---------+----------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X48:"xpc10:48" 1010 :  major_start_pcl=104   edge_private_start/end=-1/-1 exec=104 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X48:"xpc10:48"
//res2: Thread=xpc10 state=X48:"xpc10:48"
//*-------+------+---------+--------------------------------------------------------------*
//| pc    | eno  | Phaser  | Work                                                         |
//*-------+------+---------+--------------------------------------------------------------*
//| 104   | -    | R0 CTRL |                                                              |
//| 104   | 1010 | R0 DATA |                                                              |
//| 104+E | 1010 | W0 DATA | @_SINT/CC/SCALbx24_stats_lookup_probes te=te:104 scalarw(E5) |
//*-------+------+---------+--------------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X49:"xpc10:49" 1011 :  major_start_pcl=105   edge_private_start/end=-1/-1 exec=105 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X49:"xpc10:49"
//res2: Thread=xpc10 state=X49:"xpc10:49"
//*-------+------+---------+------------------------------------*
//| pc    | eno  | Phaser  | Work                               |
//*-------+------+---------+------------------------------------*
//| 105   | -    | R0 CTRL |                                    |
//| 105   | 1011 | R0 DATA |                                    |
//| 105+E | 1011 | W0 DATA | TCha3.10_V_0 te=te:105 scalarw(E6) |
//*-------+------+---------+------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X50:"xpc10:50" 1013 :  major_start_pcl=106   edge_private_start/end=107/170 exec=170 (dend=64)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X50:"xpc10:50" 1012 :  major_start_pcl=106   edge_private_start/end=-1/-1 exec=106 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X50:"xpc10:50"
//res2: Thread=xpc10 state=X50:"xpc10:50"
//*---------+------+----------+----------------------------------------------------------*
//| pc      | eno  | Phaser   | Work                                                     |
//*---------+------+----------+----------------------------------------------------------*
//| 106     | -    | R0 CTRL  |                                                          |
//| 106     | 1012 | R0 DATA  |                                                          |
//| 106+E   | 1012 | W0 DATA  | TCha3.10_V_0 te=te:106 scalarw(-TCha3.10_V_0)            |
//| 106+S   | 1013 | R0 DATA  | isMODULUS10 te=te:106 *fixed-func-ALU*(TCha3.10_V_0, E7) |
//| 107     | 1013 | R1 DATA  |                                                          |
//| 108     | 1013 | R2 DATA  |                                                          |
//| 109     | 1013 | R3 DATA  |                                                          |
//| 110     | 1013 | R4 DATA  |                                                          |
//| 111     | 1013 | R5 DATA  |                                                          |
//| 112     | 1013 | R6 DATA  |                                                          |
//| 113     | 1013 | R7 DATA  |                                                          |
//| 114     | 1013 | R8 DATA  |                                                          |
//| 115     | 1013 | R9 DATA  |                                                          |
//| 116     | 1013 | R10 DATA |                                                          |
//| 117     | 1013 | R11 DATA |                                                          |
//| 118     | 1013 | R12 DATA |                                                          |
//| 119     | 1013 | R13 DATA |                                                          |
//| 120     | 1013 | R14 DATA |                                                          |
//| 121     | 1013 | R15 DATA |                                                          |
//| 122     | 1013 | R16 DATA |                                                          |
//| 123     | 1013 | R17 DATA |                                                          |
//| 124     | 1013 | R18 DATA |                                                          |
//| 125     | 1013 | R19 DATA |                                                          |
//| 126     | 1013 | R20 DATA |                                                          |
//| 127     | 1013 | R21 DATA |                                                          |
//| 128     | 1013 | R22 DATA |                                                          |
//| 129     | 1013 | R23 DATA |                                                          |
//| 130     | 1013 | R24 DATA |                                                          |
//| 131     | 1013 | R25 DATA |                                                          |
//| 132     | 1013 | R26 DATA |                                                          |
//| 133     | 1013 | R27 DATA |                                                          |
//| 134     | 1013 | R28 DATA |                                                          |
//| 135     | 1013 | R29 DATA |                                                          |
//| 136     | 1013 | R30 DATA |                                                          |
//| 137     | 1013 | R31 DATA |                                                          |
//| 138     | 1013 | R32 DATA |                                                          |
//| 139     | 1013 | R33 DATA |                                                          |
//| 140     | 1013 | R34 DATA |                                                          |
//| 141     | 1013 | R35 DATA |                                                          |
//| 142     | 1013 | R36 DATA |                                                          |
//| 143     | 1013 | R37 DATA |                                                          |
//| 144     | 1013 | R38 DATA |                                                          |
//| 145     | 1013 | R39 DATA |                                                          |
//| 146     | 1013 | R40 DATA |                                                          |
//| 147     | 1013 | R41 DATA |                                                          |
//| 148     | 1013 | R42 DATA |                                                          |
//| 149     | 1013 | R43 DATA |                                                          |
//| 150     | 1013 | R44 DATA |                                                          |
//| 151     | 1013 | R45 DATA |                                                          |
//| 152     | 1013 | R46 DATA |                                                          |
//| 153     | 1013 | R47 DATA |                                                          |
//| 154     | 1013 | R48 DATA |                                                          |
//| 155     | 1013 | R49 DATA |                                                          |
//| 156     | 1013 | R50 DATA |                                                          |
//| 157     | 1013 | R51 DATA |                                                          |
//| 158     | 1013 | R52 DATA |                                                          |
//| 159     | 1013 | R53 DATA |                                                          |
//| 160     | 1013 | R54 DATA |                                                          |
//| 161     | 1013 | R55 DATA |                                                          |
//| 162     | 1013 | R56 DATA |                                                          |
//| 163     | 1013 | R57 DATA |                                                          |
//| 164     | 1013 | R58 DATA |                                                          |
//| 165     | 1013 | R59 DATA |                                                          |
//| 166     | 1013 | R60 DATA |                                                          |
//| 167     | 1013 | R61 DATA |                                                          |
//| 168     | 1013 | R62 DATA |                                                          |
//| 169     | 1013 | R63 DATA |                                                          |
//| 170+S   | 1013 | R64 DATA |                                                          |
//| 170+E+S | 1013 | W0 DATA  | TClo6.9_V_1 te=te:170 scalarw(E8)                        |
//*---------+------+----------+----------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X51:"xpc10:51" 1014 :  major_start_pcl=171   edge_private_start/end=172/235 exec=235 (dend=64)
//Simple greedy schedule for res2: Thread=xpc10 state=X51:"xpc10:51"
//res2: Thread=xpc10 state=X51:"xpc10:51"
//*---------+------+----------+----------------------------------------------------------*
//| pc      | eno  | Phaser   | Work                                                     |
//*---------+------+----------+----------------------------------------------------------*
//| 171     | -    | R0 CTRL  |                                                          |
//| 171+S   | 1014 | R0 DATA  | isMODULUS10 te=te:171 *fixed-func-ALU*(TCha3.10_V_0, E7) |
//| 172     | 1014 | R1 DATA  |                                                          |
//| 173     | 1014 | R2 DATA  |                                                          |
//| 174     | 1014 | R3 DATA  |                                                          |
//| 175     | 1014 | R4 DATA  |                                                          |
//| 176     | 1014 | R5 DATA  |                                                          |
//| 177     | 1014 | R6 DATA  |                                                          |
//| 178     | 1014 | R7 DATA  |                                                          |
//| 179     | 1014 | R8 DATA  |                                                          |
//| 180     | 1014 | R9 DATA  |                                                          |
//| 181     | 1014 | R10 DATA |                                                          |
//| 182     | 1014 | R11 DATA |                                                          |
//| 183     | 1014 | R12 DATA |                                                          |
//| 184     | 1014 | R13 DATA |                                                          |
//| 185     | 1014 | R14 DATA |                                                          |
//| 186     | 1014 | R15 DATA |                                                          |
//| 187     | 1014 | R16 DATA |                                                          |
//| 188     | 1014 | R17 DATA |                                                          |
//| 189     | 1014 | R18 DATA |                                                          |
//| 190     | 1014 | R19 DATA |                                                          |
//| 191     | 1014 | R20 DATA |                                                          |
//| 192     | 1014 | R21 DATA |                                                          |
//| 193     | 1014 | R22 DATA |                                                          |
//| 194     | 1014 | R23 DATA |                                                          |
//| 195     | 1014 | R24 DATA |                                                          |
//| 196     | 1014 | R25 DATA |                                                          |
//| 197     | 1014 | R26 DATA |                                                          |
//| 198     | 1014 | R27 DATA |                                                          |
//| 199     | 1014 | R28 DATA |                                                          |
//| 200     | 1014 | R29 DATA |                                                          |
//| 201     | 1014 | R30 DATA |                                                          |
//| 202     | 1014 | R31 DATA |                                                          |
//| 203     | 1014 | R32 DATA |                                                          |
//| 204     | 1014 | R33 DATA |                                                          |
//| 205     | 1014 | R34 DATA |                                                          |
//| 206     | 1014 | R35 DATA |                                                          |
//| 207     | 1014 | R36 DATA |                                                          |
//| 208     | 1014 | R37 DATA |                                                          |
//| 209     | 1014 | R38 DATA |                                                          |
//| 210     | 1014 | R39 DATA |                                                          |
//| 211     | 1014 | R40 DATA |                                                          |
//| 212     | 1014 | R41 DATA |                                                          |
//| 213     | 1014 | R42 DATA |                                                          |
//| 214     | 1014 | R43 DATA |                                                          |
//| 215     | 1014 | R44 DATA |                                                          |
//| 216     | 1014 | R45 DATA |                                                          |
//| 217     | 1014 | R46 DATA |                                                          |
//| 218     | 1014 | R47 DATA |                                                          |
//| 219     | 1014 | R48 DATA |                                                          |
//| 220     | 1014 | R49 DATA |                                                          |
//| 221     | 1014 | R50 DATA |                                                          |
//| 222     | 1014 | R51 DATA |                                                          |
//| 223     | 1014 | R52 DATA |                                                          |
//| 224     | 1014 | R53 DATA |                                                          |
//| 225     | 1014 | R54 DATA |                                                          |
//| 226     | 1014 | R55 DATA |                                                          |
//| 227     | 1014 | R56 DATA |                                                          |
//| 228     | 1014 | R57 DATA |                                                          |
//| 229     | 1014 | R58 DATA |                                                          |
//| 230     | 1014 | R59 DATA |                                                          |
//| 231     | 1014 | R60 DATA |                                                          |
//| 232     | 1014 | R61 DATA |                                                          |
//| 233     | 1014 | R62 DATA |                                                          |
//| 234     | 1014 | R63 DATA |                                                          |
//| 235+S   | 1014 | R64 DATA |                                                          |
//| 235+E+S | 1014 | W0 DATA  | TClo6.9_V_1 te=te:235 scalarw(E8)                        |
//*---------+------+----------+----------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X52:"xpc10:52" 1017 :  major_start_pcl=236   edge_private_start/end=-1/-1 exec=237 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X52:"xpc10:52" 1016 :  major_start_pcl=236   edge_private_start/end=-1/-1 exec=237 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X52:"xpc10:52" 1015 :  major_start_pcl=236   edge_private_start/end=-1/-1 exec=237 (dend=1)
//Simple greedy schedule for res2: Thread=xpc10 state=X52:"xpc10:52"
//res2: Thread=xpc10 state=X52:"xpc10:52"
//*-------+------+---------+----------------------------------------------------------------------------------------------------------------------------------------------------*
//| pc    | eno  | Phaser  | Work                                                                                                                                               |
//*-------+------+---------+----------------------------------------------------------------------------------------------------------------------------------------------------*
//| 236   | -    | R0 CTRL | @_SINT/CC/MAPR10NoCE3_ARA0 te=te:236 read(TClo6.9_V_1) @_SINT/CC/MAPR10NoCE2_ARA0 te=te:236 read(TClo6.9_V_1) @_SINT/CC/MAPR10NoCE1_ARA0 te=te:23\ |
//|       |      |         | 6 read(TClo6.9_V_1) @_SINT/CC/MAPR10NoCE0_ARA0 te=te:236 read(TClo6.9_V_1)                                                                         |
//| 237   | -    | R1 CTRL |                                                                                                                                                    |
//| 236   | 1015 | R0 DATA |                                                                                                                                                    |
//| 237   | 1015 | R1 DATA |                                                                                                                                                    |
//| 237+E | 1015 | W0 DATA | TCl6._SPILL_256 te=te:237 scalarw(-5) TTMT4Main_V_14 te=te:237 scalarw(S32'-5I)                                                                    |
//| 236   | 1016 | R0 DATA | @_SINT/CC/MAPR12NoCE3_ARB0 te=te:236 read(TClo6.9_V_1) @_SINT/CC/MAPR12NoCE2_ARB0 te=te:236 read(TClo6.9_V_1) @_SINT/CC/MAPR12NoCE1_ARB0 te=te:23\ |
//|       |      |         | 6 read(TClo6.9_V_1) @_SINT/CC/MAPR12NoCE0_ARB0 te=te:236 read(TClo6.9_V_1)                                                                         |
//| 237   | 1016 | R1 DATA |                                                                                                                                                    |
//| 237+E | 1016 | W0 DATA | TClo6.9_V_2 te=te:237 scalarw(E9)                                                                                                                  |
//| 236   | 1017 | R0 DATA |                                                                                                                                                    |
//| 237   | 1017 | R1 DATA |                                                                                                                                                    |
//| 237+E | 1017 | W0 DATA | TClo6.9_V_0 te=te:237 scalarw(1+TClo6.9_V_0)                                                                                                       |
//*-------+------+---------+----------------------------------------------------------------------------------------------------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X53:"xpc10:53" 1020 :  major_start_pcl=238   edge_private_start/end=-1/-1 exec=238 (dend=0)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X53:"xpc10:53" 1019 :  major_start_pcl=238   edge_private_start/end=-1/-1 exec=238 (dend=0)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X53:"xpc10:53" 1018 :  major_start_pcl=238   edge_private_start/end=-1/-1 exec=238 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X53:"xpc10:53"
//res2: Thread=xpc10 state=X53:"xpc10:53"
//*-------+------+---------+--------------------------------------------------*
//| pc    | eno  | Phaser  | Work                                             |
//*-------+------+---------+--------------------------------------------------*
//| 238   | -    | R0 CTRL |                                                  |
//| 238   | 1018 | R0 DATA |                                                  |
//| 238+E | 1018 | W0 DATA | TTMT4Main_V_9 te=te:238 scalarw(1+TTMT4Main_V_9) |
//| 238   | 1019 | R0 DATA |                                                  |
//| 238+E | 1019 | W0 DATA | TTMT4Main_V_8 te=te:238 scalarw(1+TTMT4Main_V_8) |
//| 238   | 1020 | R0 DATA |                                                  |
//| 238+E | 1020 | W0 DATA | TTMT4Main_V_8 te=te:238 scalarw(1+TTMT4Main_V_8) |
//*-------+------+---------+--------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X54:"xpc10:54" 1021 :  major_start_pcl=239   edge_private_start/end=240/240 exec=240 (dend=1)
//Simple greedy schedule for res2: Thread=xpc10 state=X54:"xpc10:54"
//res2: Thread=xpc10 state=X54:"xpc10:54"
//*-------+------+---------+-----------------------------------------------------*
//| pc    | eno  | Phaser  | Work                                                |
//*-------+------+---------+-----------------------------------------------------*
//| 239   | -    | R0 CTRL |                                                     |
//| 239   | 1021 | R0 DATA | @64_US/CC/SCALbx26_ARA0 te=te:239 read(TClo6.9_V_2) |
//| 240   | 1021 | R1 DATA |                                                     |
//| 240+E | 1021 | W0 DATA | TTMT4Main_V_13 te=te:240 scalarw(E10)               |
//*-------+------+---------+-----------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X55:"xpc10:55" 1022 :  major_start_pcl=241   edge_private_start/end=-1/-1 exec=241 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X55:"xpc10:55"
//res2: Thread=xpc10 state=X55:"xpc10:55"
//*-------+------+---------+-------------------------------------------------------------------------------*
//| pc    | eno  | Phaser  | Work                                                                          |
//*-------+------+---------+-------------------------------------------------------------------------------*
//| 241   | -    | R0 CTRL |                                                                               |
//| 241   | 1022 | R0 DATA |                                                                               |
//| 241+E | 1022 | W0 DATA | TCl6._SPILL_256 te=te:241 scalarw(0) TTMT4Main_V_14 te=te:241 scalarw(S32'0I) |
//*-------+------+---------+-------------------------------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X56:"xpc10:56" 1025 :  major_start_pcl=242   edge_private_start/end=-1/-1 exec=242 (dend=0)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X56:"xpc10:56" 1024 :  major_start_pcl=242   edge_private_start/end=243/243 exec=243 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X56:"xpc10:56" 1023 :  major_start_pcl=242   edge_private_start/end=-1/-1 exec=242 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X56:"xpc10:56"
//res2: Thread=xpc10 state=X56:"xpc10:56"
//*-------+------+---------+----------------------------------------------------------------------------------------------------------------------------------------------------*
//| pc    | eno  | Phaser  | Work                                                                                                                                               |
//*-------+------+---------+----------------------------------------------------------------------------------------------------------------------------------------------------*
//| 242   | -    | R0 CTRL |                                                                                                                                                    |
//| 242   | 1023 | R0 DATA |                                                                                                                                                    |
//| 242+E | 1023 | W0 DATA | TCl6._SPILL_256 te=te:242 scalarw(-5) TTMT4Main_V_14 te=te:242 scalarw(S32'-5I) @_SINT/CC/SCALbx24_stats_lookup_probes te=te:242 scalarw(E5)       |
//| 242   | 1024 | R0 DATA | @_SINT/CC/MAPR12NoCE3_ARB0 te=te:242 read(TClo6.9_V_1) @_SINT/CC/MAPR12NoCE2_ARB0 te=te:242 read(TClo6.9_V_1) @_SINT/CC/MAPR12NoCE1_ARB0 te=te:24\ |
//|       |      |         | 2 read(TClo6.9_V_1) @_SINT/CC/MAPR12NoCE0_ARB0 te=te:242 read(TClo6.9_V_1)                                                                         |
//| 243   | 1024 | R1 DATA |                                                                                                                                                    |
//| 243+E | 1024 | W0 DATA | TClo6.9_V_2 te=te:243 scalarw(E9)                                                                                                                  |
//| 242   | 1025 | R0 DATA |                                                                                                                                                    |
//| 242+E | 1025 | W0 DATA | TCl6._SPILL_256 te=te:242 scalarw(-5) TTMT4Main_V_14 te=te:242 scalarw(S32'-5I) @_SINT/CC/SCALbx24_stats_lookup_probes te=te:242 scalarw(E5)       |
//*-------+------+---------+----------------------------------------------------------------------------------------------------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X57:"xpc10:57" 1026 :  major_start_pcl=244   edge_private_start/end=-1/-1 exec=244 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X57:"xpc10:57"
//res2: Thread=xpc10 state=X57:"xpc10:57"
//*-------+------+---------+-------------------------------------*
//| pc    | eno  | Phaser  | Work                                |
//*-------+------+---------+-------------------------------------*
//| 244   | -    | R0 CTRL |                                     |
//| 244   | 1026 | R0 DATA |                                     |
//| 244+E | 1026 | W0 DATA | TTMT4Main_V_5 te=te:244 scalarw(E2) |
//*-------+------+---------+-------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X58:"xpc10:58" 1027 :  major_start_pcl=245   edge_private_start/end=-1/-1 exec=245 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X58:"xpc10:58"
//res2: Thread=xpc10 state=X58:"xpc10:58"
//*-------+------+---------+------------------------------------------------------------------------*
//| pc    | eno  | Phaser  | Work                                                                   |
//*-------+------+---------+------------------------------------------------------------------------*
//| 245   | -    | R0 CTRL |                                                                        |
//| 245   | 1027 | R0 DATA |                                                                        |
//| 245+E | 1027 | W0 DATA | TDGe1.4_V_0 te=te:245 scalarw(E3) fastspilldup12 te=te:245 scalarw(E3) |
//*-------+------+---------+------------------------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X59:"xpc10:59" 1028 :  major_start_pcl=246   edge_private_start/end=-1/-1 exec=246 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X59:"xpc10:59"
//res2: Thread=xpc10 state=X59:"xpc10:59"
//*-------+------+---------+----------------------------------------------------------------*
//| pc    | eno  | Phaser  | Work                                                           |
//*-------+------+---------+----------------------------------------------------------------*
//| 246   | -    | R0 CTRL |                                                                |
//| 246   | 1028 | R0 DATA |                                                                |
//| 246+E | 1028 | W0 DATA | @64_US/CC/SCALbx28_dk te=te:246 scalarw(S64'1I+fastspilldup12) |
//*-------+------+---------+----------------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X60:"xpc10:60" 1029 :  major_start_pcl=247   edge_private_start/end=-1/-1 exec=247 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X60:"xpc10:60"
//res2: Thread=xpc10 state=X60:"xpc10:60"
//*-------+------+---------+----------------------------------------------------------------------------------------------------*
//| pc    | eno  | Phaser  | Work                                                                                               |
//*-------+------+---------+----------------------------------------------------------------------------------------------------*
//| 247   | -    | R0 CTRL |                                                                                                    |
//| 247   | 1029 | R0 DATA |                                                                                                    |
//| 247+E | 1029 | W0 DATA | TCin1.9_V_0 te=te:247 scalarw(C(TTMT4Main_V_5)) TTMT4Main_V_6 te=te:247 scalarw(C64u(TDGe1.4_V_0)) |
//*-------+------+---------+----------------------------------------------------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X61:"xpc10:61" 1030 :  major_start_pcl=248   edge_private_start/end=-1/-1 exec=248 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X61:"xpc10:61"
//res2: Thread=xpc10 state=X61:"xpc10:61"
//*-------+------+---------+-------------------------------------------------------------------*
//| pc    | eno  | Phaser  | Work                                                              |
//*-------+------+---------+-------------------------------------------------------------------*
//| 248   | -    | R0 CTRL |                                                                   |
//| 248   | 1030 | R0 DATA |                                                                   |
//| 248+E | 1030 | W0 DATA | TCin1.9_V_2 te=te:248 scalarw(0) TCin1.9_V_1 te=te:248 scalarw(0) |
//*-------+------+---------+-------------------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X62:"xpc10:62" 1033 :  major_start_pcl=249   edge_private_start/end=-1/-1 exec=249 (dend=0)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X62:"xpc10:62" 1032 :  major_start_pcl=249   edge_private_start/end=-1/-1 exec=249 (dend=0)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X62:"xpc10:62" 1031 :  major_start_pcl=249   edge_private_start/end=-1/-1 exec=249 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X62:"xpc10:62"
//res2: Thread=xpc10 state=X62:"xpc10:62"
//*-------+------+---------+--------------------------------------------------------------------------------*
//| pc    | eno  | Phaser  | Work                                                                           |
//*-------+------+---------+--------------------------------------------------------------------------------*
//| 249   | -    | R0 CTRL |                                                                                |
//| 249   | 1031 | R0 DATA |                                                                                |
//| 249+E | 1031 | W0 DATA | TTMT4Main_V_7 te=te:249 scalarw(S32'-4I) TCi1._SPILL_256 te=te:249 scalarw(-4) |
//| 249   | 1032 | R0 DATA |                                                                                |
//| 249+E | 1032 | W0 DATA | TTMT4Main_V_7 te=te:249 scalarw(S32'-2I) TCi1._SPILL_256 te=te:249 scalarw(-2) |
//| 249   | 1033 | R0 DATA |                                                                                |
//| 249+E | 1033 | W0 DATA | fastspilldup16 te=te:249 scalarw(E11)                                          |
//*-------+------+---------+--------------------------------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X63:"xpc10:63" 1035 :  major_start_pcl=250   edge_private_start/end=-1/-1 exec=250 (dend=0)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X63:"xpc10:63" 1034 :  major_start_pcl=250   edge_private_start/end=-1/-1 exec=250 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X63:"xpc10:63"
//res2: Thread=xpc10 state=X63:"xpc10:63"
//*-------+------+---------+--------------------------------------------------*
//| pc    | eno  | Phaser  | Work                                             |
//*-------+------+---------+--------------------------------------------------*
//| 250   | -    | R0 CTRL |                                                  |
//| 250   | 1034 | R0 DATA |                                                  |
//| 250+E | 1034 | W0 DATA | TTMT4Main_V_3 te=te:250 scalarw(1+TTMT4Main_V_3) |
//| 250   | 1035 | R0 DATA |                                                  |
//| 250+E | 1035 | W0 DATA | TTMT4Main_V_2 te=te:250 scalarw(1+TTMT4Main_V_2) |
//*-------+------+---------+--------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X64:"xpc10:64" 1036 :  major_start_pcl=251   edge_private_start/end=-1/-1 exec=251 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X64:"xpc10:64"
//res2: Thread=xpc10 state=X64:"xpc10:64"
//*-------+------+---------+--------------------------------------------------*
//| pc    | eno  | Phaser  | Work                                             |
//*-------+------+---------+--------------------------------------------------*
//| 251   | -    | R0 CTRL |                                                  |
//| 251   | 1036 | R0 DATA |                                                  |
//| 251+E | 1036 | W0 DATA | TTMT4Main_V_2 te=te:251 scalarw(1+TTMT4Main_V_2) |
//*-------+------+---------+--------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X65:"xpc10:65" 1037 :  major_start_pcl=252   edge_private_start/end=-1/-1 exec=252 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X65:"xpc10:65"
//res2: Thread=xpc10 state=X65:"xpc10:65"
//*-------+------+---------+--------------------------------------------------*
//| pc    | eno  | Phaser  | Work                                             |
//*-------+------+---------+--------------------------------------------------*
//| 252   | -    | R0 CTRL |                                                  |
//| 252   | 1037 | R0 DATA |                                                  |
//| 252+E | 1037 | W0 DATA | TTMT4Main_V_4 te=te:252 scalarw(1+TTMT4Main_V_4) |
//*-------+------+---------+--------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X66:"xpc10:66" 1039 :  major_start_pcl=253   edge_private_start/end=-1/-1 exec=253 (dend=0)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X66:"xpc10:66" 1038 :  major_start_pcl=253   edge_private_start/end=-1/-1 exec=253 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X66:"xpc10:66"
//res2: Thread=xpc10 state=X66:"xpc10:66"
//*-------+------+---------+------------------------------------------------*
//| pc    | eno  | Phaser  | Work                                           |
//*-------+------+---------+------------------------------------------------*
//| 253   | -    | R0 CTRL |                                                |
//| 253   | 1038 | R0 DATA |                                                |
//| 253+E | 1038 | W0 DATA |  W/P:Data Entered  PLI:Cuckoo cache inserte... |
//| 253   | 1039 | R0 DATA |                                                |
//| 253+E | 1039 | W0 DATA | @_SINT/CC/SCALbx28_seed te=te:253 scalarw(E1)  |
//*-------+------+---------+------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X67:"xpc10:67" 1040 :  major_start_pcl=254   edge_private_start/end=-1/-1 exec=254 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X67:"xpc10:67"
//res2: Thread=xpc10 state=X67:"xpc10:67"
//*-------+------+---------+-------------------------------------------------------------------------------------------------------------------*
//| pc    | eno  | Phaser  | Work                                                                                                              |
//*-------+------+---------+-------------------------------------------------------------------------------------------------------------------*
//| 254   | -    | R0 CTRL |                                                                                                                   |
//| 254   | 1040 | R0 DATA |                                                                                                                   |
//| 254+E | 1040 | W0 DATA | @_SINT/CC/SCALbx24_next_free te=te:254 scalarw(1+fastspilldup16) TCin1.9_V_3 te=te:254 scalarw(C(fastspilldup16)) |
//*-------+------+---------+-------------------------------------------------------------------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X68:"xpc10:68" 1041 :  major_start_pcl=255   edge_private_start/end=256/256 exec=255 (dend=1)
//Simple greedy schedule for res2: Thread=xpc10 state=X68:"xpc10:68"
//res2: Thread=xpc10 state=X68:"xpc10:68"
//*-------+------+---------+----------------------------------------------------------------------------------------------------------------------------*
//| pc    | eno  | Phaser  | Work                                                                                                                       |
//*-------+------+---------+----------------------------------------------------------------------------------------------------------------------------*
//| 255   | -    | R0 CTRL |                                                                                                                            |
//| 255   | 1041 | R0 DATA |                                                                                                                            |
//| 255+E | 1041 | W0 DATA | @64_US/CC/SCALbx26_ARA0 te=te:255 write(C(TCin1.9_V_3), C64u(TTMT4Main_V_6)) TCin1.9_V_2 te=te:255 scalarw(C(TCin1.9_V_3)) |
//| 256   | 1041 | W1 DATA |                                                                                                                            |
//*-------+------+---------+----------------------------------------------------------------------------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X69:"xpc10:69" 1042 :  major_start_pcl=257   edge_private_start/end=-1/-1 exec=257 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X69:"xpc10:69"
//res2: Thread=xpc10 state=X69:"xpc10:69"
//*-------+------+---------+---------------------------------------------------------*
//| pc    | eno  | Phaser  | Work                                                    |
//*-------+------+---------+---------------------------------------------------------*
//| 257   | -    | R0 CTRL |                                                         |
//| 257   | 1042 | R0 DATA |                                                         |
//| 257+E | 1042 | W0 DATA | @_SINT/CC/SCALbx24_stats_inserts te=te:257 scalarw(E12) |
//*-------+------+---------+---------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X70:"xpc10:70" 1043 :  major_start_pcl=258   edge_private_start/end=-1/-1 exec=258 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X70:"xpc10:70"
//res2: Thread=xpc10 state=X70:"xpc10:70"
//*-------+------+---------+-------------------------------------------------------------------*
//| pc    | eno  | Phaser  | Work                                                              |
//*-------+------+---------+-------------------------------------------------------------------*
//| 258   | -    | R0 CTRL |                                                                   |
//| 258   | 1043 | R0 DATA |                                                                   |
//| 258+E | 1043 | W0 DATA | TCin1.9_V_4 te=te:258 scalarw(0) TCin1.9_V_5 te=te:258 scalarw(0) |
//*-------+------+---------+-------------------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X71:"xpc10:71" 1070 :  major_start_pcl=259   edge_private_start/end=-1/-1 exec=259 (dend=0)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X71:"xpc10:71" 1069 :  major_start_pcl=259   edge_private_start/end=-1/-1 exec=259 (dend=0)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X71:"xpc10:71" 1068 :  major_start_pcl=259   edge_private_start/end=283/283 exec=259 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X71:"xpc10:71" 1067 :  major_start_pcl=259   edge_private_start/end=282/282 exec=259 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X71:"xpc10:71" 1066 :  major_start_pcl=259   edge_private_start/end=281/281 exec=259 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X71:"xpc10:71" 1065 :  major_start_pcl=259   edge_private_start/end=280/280 exec=259 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X71:"xpc10:71" 1064 :  major_start_pcl=259   edge_private_start/end=279/279 exec=259 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X71:"xpc10:71" 1063 :  major_start_pcl=259   edge_private_start/end=278/278 exec=259 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X71:"xpc10:71" 1062 :  major_start_pcl=259   edge_private_start/end=277/277 exec=259 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X71:"xpc10:71" 1061 :  major_start_pcl=259   edge_private_start/end=276/276 exec=259 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X71:"xpc10:71" 1060 :  major_start_pcl=259   edge_private_start/end=275/275 exec=259 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X71:"xpc10:71" 1059 :  major_start_pcl=259   edge_private_start/end=274/274 exec=259 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X71:"xpc10:71" 1058 :  major_start_pcl=259   edge_private_start/end=273/273 exec=259 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X71:"xpc10:71" 1057 :  major_start_pcl=259   edge_private_start/end=272/272 exec=259 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X71:"xpc10:71" 1056 :  major_start_pcl=259   edge_private_start/end=271/271 exec=259 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X71:"xpc10:71" 1055 :  major_start_pcl=259   edge_private_start/end=270/270 exec=259 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X71:"xpc10:71" 1054 :  major_start_pcl=259   edge_private_start/end=269/269 exec=259 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X71:"xpc10:71" 1053 :  major_start_pcl=259   edge_private_start/end=268/268 exec=259 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X71:"xpc10:71" 1052 :  major_start_pcl=259   edge_private_start/end=267/267 exec=259 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X71:"xpc10:71" 1051 :  major_start_pcl=259   edge_private_start/end=266/266 exec=259 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X71:"xpc10:71" 1050 :  major_start_pcl=259   edge_private_start/end=265/265 exec=259 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X71:"xpc10:71" 1049 :  major_start_pcl=259   edge_private_start/end=264/264 exec=259 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X71:"xpc10:71" 1048 :  major_start_pcl=259   edge_private_start/end=263/263 exec=259 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X71:"xpc10:71" 1047 :  major_start_pcl=259   edge_private_start/end=262/262 exec=259 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X71:"xpc10:71" 1046 :  major_start_pcl=259   edge_private_start/end=261/261 exec=259 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X71:"xpc10:71" 1045 :  major_start_pcl=259   edge_private_start/end=260/260 exec=259 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X71:"xpc10:71" 1044 :  major_start_pcl=259   edge_private_start/end=-1/-1 exec=259 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X71:"xpc10:71"
//res2: Thread=xpc10 state=X71:"xpc10:71"
//*-------+------+---------+-------------------------------------------------------------------------------------------------------------------------------------------------*
//| pc    | eno  | Phaser  | Work                                                                                                                                            |
//*-------+------+---------+-------------------------------------------------------------------------------------------------------------------------------------------------*
//| 259   | -    | R0 CTRL |                                                                                                                                                 |
//| 259   | 1044 | R0 DATA |                                                                                                                                                 |
//| 259+E | 1044 | W0 DATA | TCin1.9_V_1 te=te:259 scalarw(1+TCin1.9_V_1) @_SINT/CC/SCALbx24_stats_insert_probes te=te:259 scalarw(E13)  PLI:Eviction %u needed              |
//| 259   | 1045 | R0 DATA |                                                                                                                                                 |
//| 259+E | 1045 | W0 DATA | @_SINT/CC/MAPR10NoCE3_ARA0 te=te:259 write(TCin1.9_V_5, C(TCin1.9_V_0)) @_SINT/CC/MAPR12NoCE3_ARB0 te=te:259 write(TCin1.9_V_5, C(TCin1.9_V_2)) |
//| 260   | 1045 | W1 DATA |                                                                                                                                                 |
//| 259   | 1046 | R0 DATA |                                                                                                                                                 |
//| 259+E | 1046 | W0 DATA | @_SINT/CC/MAPR10NoCE3_ARA0 te=te:259 write(TCin1.9_V_5, C(TCin1.9_V_0)) @_SINT/CC/MAPR12NoCE2_ARB0 te=te:259 write(TCin1.9_V_5, C(TCin1.9_V_2)) |
//| 261   | 1046 | W1 DATA |                                                                                                                                                 |
//| 259   | 1047 | R0 DATA |                                                                                                                                                 |
//| 259+E | 1047 | W0 DATA | @_SINT/CC/MAPR10NoCE3_ARA0 te=te:259 write(TCin1.9_V_5, C(TCin1.9_V_0)) @_SINT/CC/MAPR12NoCE1_ARB0 te=te:259 write(TCin1.9_V_5, C(TCin1.9_V_2)) |
//| 262   | 1047 | W1 DATA |                                                                                                                                                 |
//| 259   | 1048 | R0 DATA |                                                                                                                                                 |
//| 259+E | 1048 | W0 DATA | @_SINT/CC/MAPR10NoCE3_ARA0 te=te:259 write(TCin1.9_V_5, C(TCin1.9_V_0)) @_SINT/CC/MAPR12NoCE0_ARB0 te=te:259 write(TCin1.9_V_5, C(TCin1.9_V_2)) |
//| 263   | 1048 | W1 DATA |                                                                                                                                                 |
//| 259   | 1049 | R0 DATA |                                                                                                                                                 |
//| 259+E | 1049 | W0 DATA | @_SINT/CC/MAPR10NoCE3_ARA0 te=te:259 write(TCin1.9_V_5, C(TCin1.9_V_0)) TCi1._SPILL_256 te=te:259 scalarw(0)                                    |
//| 264   | 1049 | W1 DATA |                                                                                                                                                 |
//| 259   | 1050 | R0 DATA |                                                                                                                                                 |
//| 259+E | 1050 | W0 DATA | @_SINT/CC/MAPR10NoCE2_ARA0 te=te:259 write(TCin1.9_V_5, C(TCin1.9_V_0)) @_SINT/CC/MAPR12NoCE3_ARB0 te=te:259 write(TCin1.9_V_5, C(TCin1.9_V_2)) |
//| 265   | 1050 | W1 DATA |                                                                                                                                                 |
//| 259   | 1051 | R0 DATA |                                                                                                                                                 |
//| 259+E | 1051 | W0 DATA | @_SINT/CC/MAPR10NoCE2_ARA0 te=te:259 write(TCin1.9_V_5, C(TCin1.9_V_0)) @_SINT/CC/MAPR12NoCE2_ARB0 te=te:259 write(TCin1.9_V_5, C(TCin1.9_V_2)) |
//| 266   | 1051 | W1 DATA |                                                                                                                                                 |
//| 259   | 1052 | R0 DATA |                                                                                                                                                 |
//| 259+E | 1052 | W0 DATA | @_SINT/CC/MAPR10NoCE2_ARA0 te=te:259 write(TCin1.9_V_5, C(TCin1.9_V_0)) @_SINT/CC/MAPR12NoCE1_ARB0 te=te:259 write(TCin1.9_V_5, C(TCin1.9_V_2)) |
//| 267   | 1052 | W1 DATA |                                                                                                                                                 |
//| 259   | 1053 | R0 DATA |                                                                                                                                                 |
//| 259+E | 1053 | W0 DATA | @_SINT/CC/MAPR10NoCE2_ARA0 te=te:259 write(TCin1.9_V_5, C(TCin1.9_V_0)) @_SINT/CC/MAPR12NoCE0_ARB0 te=te:259 write(TCin1.9_V_5, C(TCin1.9_V_2)) |
//| 268   | 1053 | W1 DATA |                                                                                                                                                 |
//| 259   | 1054 | R0 DATA |                                                                                                                                                 |
//| 259+E | 1054 | W0 DATA | @_SINT/CC/MAPR10NoCE2_ARA0 te=te:259 write(TCin1.9_V_5, C(TCin1.9_V_0)) TCi1._SPILL_256 te=te:259 scalarw(0)                                    |
//| 269   | 1054 | W1 DATA |                                                                                                                                                 |
//| 259   | 1055 | R0 DATA |                                                                                                                                                 |
//| 259+E | 1055 | W0 DATA | @_SINT/CC/MAPR10NoCE1_ARA0 te=te:259 write(TCin1.9_V_5, C(TCin1.9_V_0)) @_SINT/CC/MAPR12NoCE3_ARB0 te=te:259 write(TCin1.9_V_5, C(TCin1.9_V_2)) |
//| 270   | 1055 | W1 DATA |                                                                                                                                                 |
//| 259   | 1056 | R0 DATA |                                                                                                                                                 |
//| 259+E | 1056 | W0 DATA | @_SINT/CC/MAPR10NoCE1_ARA0 te=te:259 write(TCin1.9_V_5, C(TCin1.9_V_0)) @_SINT/CC/MAPR12NoCE2_ARB0 te=te:259 write(TCin1.9_V_5, C(TCin1.9_V_2)) |
//| 271   | 1056 | W1 DATA |                                                                                                                                                 |
//| 259   | 1057 | R0 DATA |                                                                                                                                                 |
//| 259+E | 1057 | W0 DATA | @_SINT/CC/MAPR10NoCE1_ARA0 te=te:259 write(TCin1.9_V_5, C(TCin1.9_V_0)) @_SINT/CC/MAPR12NoCE1_ARB0 te=te:259 write(TCin1.9_V_5, C(TCin1.9_V_2)) |
//| 272   | 1057 | W1 DATA |                                                                                                                                                 |
//| 259   | 1058 | R0 DATA |                                                                                                                                                 |
//| 259+E | 1058 | W0 DATA | @_SINT/CC/MAPR10NoCE1_ARA0 te=te:259 write(TCin1.9_V_5, C(TCin1.9_V_0)) @_SINT/CC/MAPR12NoCE0_ARB0 te=te:259 write(TCin1.9_V_5, C(TCin1.9_V_2)) |
//| 273   | 1058 | W1 DATA |                                                                                                                                                 |
//| 259   | 1059 | R0 DATA |                                                                                                                                                 |
//| 259+E | 1059 | W0 DATA | @_SINT/CC/MAPR10NoCE1_ARA0 te=te:259 write(TCin1.9_V_5, C(TCin1.9_V_0)) TCi1._SPILL_256 te=te:259 scalarw(0)                                    |
//| 274   | 1059 | W1 DATA |                                                                                                                                                 |
//| 259   | 1060 | R0 DATA |                                                                                                                                                 |
//| 259+E | 1060 | W0 DATA | @_SINT/CC/MAPR10NoCE0_ARA0 te=te:259 write(TCin1.9_V_5, C(TCin1.9_V_0)) @_SINT/CC/MAPR12NoCE3_ARB0 te=te:259 write(TCin1.9_V_5, C(TCin1.9_V_2)) |
//| 275   | 1060 | W1 DATA |                                                                                                                                                 |
//| 259   | 1061 | R0 DATA |                                                                                                                                                 |
//| 259+E | 1061 | W0 DATA | @_SINT/CC/MAPR10NoCE0_ARA0 te=te:259 write(TCin1.9_V_5, C(TCin1.9_V_0)) @_SINT/CC/MAPR12NoCE2_ARB0 te=te:259 write(TCin1.9_V_5, C(TCin1.9_V_2)) |
//| 276   | 1061 | W1 DATA |                                                                                                                                                 |
//| 259   | 1062 | R0 DATA |                                                                                                                                                 |
//| 259+E | 1062 | W0 DATA | @_SINT/CC/MAPR10NoCE0_ARA0 te=te:259 write(TCin1.9_V_5, C(TCin1.9_V_0)) @_SINT/CC/MAPR12NoCE1_ARB0 te=te:259 write(TCin1.9_V_5, C(TCin1.9_V_2)) |
//| 277   | 1062 | W1 DATA |                                                                                                                                                 |
//| 259   | 1063 | R0 DATA |                                                                                                                                                 |
//| 259+E | 1063 | W0 DATA | @_SINT/CC/MAPR10NoCE0_ARA0 te=te:259 write(TCin1.9_V_5, C(TCin1.9_V_0)) @_SINT/CC/MAPR12NoCE0_ARB0 te=te:259 write(TCin1.9_V_5, C(TCin1.9_V_2)) |
//| 278   | 1063 | W1 DATA |                                                                                                                                                 |
//| 259   | 1064 | R0 DATA |                                                                                                                                                 |
//| 259+E | 1064 | W0 DATA | @_SINT/CC/MAPR10NoCE0_ARA0 te=te:259 write(TCin1.9_V_5, C(TCin1.9_V_0)) TCi1._SPILL_256 te=te:259 scalarw(0)                                    |
//| 279   | 1064 | W1 DATA |                                                                                                                                                 |
//| 259   | 1065 | R0 DATA |                                                                                                                                                 |
//| 259+E | 1065 | W0 DATA | @_SINT/CC/MAPR12NoCE3_ARB0 te=te:259 write(TCin1.9_V_5, C(TCin1.9_V_2)) TCi1._SPILL_256 te=te:259 scalarw(0)                                    |
//| 280   | 1065 | W1 DATA |                                                                                                                                                 |
//| 259   | 1066 | R0 DATA |                                                                                                                                                 |
//| 259+E | 1066 | W0 DATA | @_SINT/CC/MAPR12NoCE2_ARB0 te=te:259 write(TCin1.9_V_5, C(TCin1.9_V_2)) TCi1._SPILL_256 te=te:259 scalarw(0)                                    |
//| 281   | 1066 | W1 DATA |                                                                                                                                                 |
//| 259   | 1067 | R0 DATA |                                                                                                                                                 |
//| 259+E | 1067 | W0 DATA | @_SINT/CC/MAPR12NoCE1_ARB0 te=te:259 write(TCin1.9_V_5, C(TCin1.9_V_2)) TCi1._SPILL_256 te=te:259 scalarw(0)                                    |
//| 282   | 1067 | W1 DATA |                                                                                                                                                 |
//| 259   | 1068 | R0 DATA |                                                                                                                                                 |
//| 259+E | 1068 | W0 DATA | @_SINT/CC/MAPR12NoCE0_ARB0 te=te:259 write(TCin1.9_V_5, C(TCin1.9_V_2)) TCi1._SPILL_256 te=te:259 scalarw(0)                                    |
//| 283   | 1068 | W1 DATA |                                                                                                                                                 |
//| 259   | 1069 | R0 DATA |                                                                                                                                                 |
//| 259+E | 1069 | W0 DATA | TTMT4Main_V_7 te=te:259 scalarw(S32'0I) TCi1._SPILL_256 te=te:259 scalarw(0)                                                                    |
//| 259   | 1070 | R0 DATA |                                                                                                                                                 |
//| 259+E | 1070 | W0 DATA | TCin1.9_V_1 te=te:259 scalarw(1+TCin1.9_V_1) @_SINT/CC/SCALbx24_stats_insert_probes te=te:259 scalarw(E13)  PLI:Eviction %u needed              |
//*-------+------+---------+-------------------------------------------------------------------------------------------------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X72:"xpc10:72" 1071 :  major_start_pcl=284   edge_private_start/end=-1/-1 exec=284 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X72:"xpc10:72"
//res2: Thread=xpc10 state=X72:"xpc10:72"
//*-------+------+---------+------------------------------------------------------------------*
//| pc    | eno  | Phaser  | Work                                                             |
//*-------+------+---------+------------------------------------------------------------------*
//| 284   | -    | R0 CTRL |                                                                  |
//| 284   | 1071 | R0 DATA |                                                                  |
//| 284+E | 1071 | W0 DATA | @_SINT/CC/SCALbx24_stats_insert_evictions te=te:284 scalarw(E14) |
//*-------+------+---------+------------------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X73:"xpc10:73" 1072 :  major_start_pcl=285   edge_private_start/end=286/286 exec=286 (dend=1)
//Simple greedy schedule for res2: Thread=xpc10 state=X73:"xpc10:73"
//res2: Thread=xpc10 state=X73:"xpc10:73"
//*-------+------+---------+----------------------------------------------------------------------------------------------------------------------------------------------------*
//| pc    | eno  | Phaser  | Work                                                                                                                                               |
//*-------+------+---------+----------------------------------------------------------------------------------------------------------------------------------------------------*
//| 285   | -    | R0 CTRL |                                                                                                                                                    |
//| 285   | 1072 | R0 DATA | @_SINT/CC/MAPR10NoCE3_ARA0 te=te:285 read(TCin1.9_V_5) @_SINT/CC/MAPR10NoCE2_ARA0 te=te:285 read(TCin1.9_V_5) @_SINT/CC/MAPR10NoCE1_ARA0 te=te:28\ |
//|       |      |         | 5 read(TCin1.9_V_5) @_SINT/CC/MAPR10NoCE0_ARA0 te=te:285 read(TCin1.9_V_5)                                                                         |
//| 286   | 1072 | R1 DATA |                                                                                                                                                    |
//| 286+E | 1072 | W0 DATA | TCin1.9_V_6 te=te:286 scalarw(E15)                                                                                                                 |
//*-------+------+---------+----------------------------------------------------------------------------------------------------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X74:"xpc10:74" 1073 :  major_start_pcl=287   edge_private_start/end=288/288 exec=288 (dend=1)
//Simple greedy schedule for res2: Thread=xpc10 state=X74:"xpc10:74"
//res2: Thread=xpc10 state=X74:"xpc10:74"
//*-------+------+---------+----------------------------------------------------------------------------------------------------------------------------------------------------*
//| pc    | eno  | Phaser  | Work                                                                                                                                               |
//*-------+------+---------+----------------------------------------------------------------------------------------------------------------------------------------------------*
//| 287   | -    | R0 CTRL |                                                                                                                                                    |
//| 287   | 1073 | R0 DATA | @_SINT/CC/MAPR12NoCE3_ARB0 te=te:287 read(TCin1.9_V_5) @_SINT/CC/MAPR12NoCE2_ARB0 te=te:287 read(TCin1.9_V_5) @_SINT/CC/MAPR12NoCE1_ARB0 te=te:28\ |
//|       |      |         | 7 read(TCin1.9_V_5) @_SINT/CC/MAPR12NoCE0_ARB0 te=te:287 read(TCin1.9_V_5)                                                                         |
//| 288   | 1073 | R1 DATA |                                                                                                                                                    |
//| 288+E | 1073 | W0 DATA | TCin1.9_V_7 te=te:288 scalarw(E16)                                                                                                                 |
//*-------+------+---------+----------------------------------------------------------------------------------------------------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X75:"xpc10:75" 1098 :  major_start_pcl=289   edge_private_start/end=-1/-1 exec=289 (dend=0)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X75:"xpc10:75" 1097 :  major_start_pcl=289   edge_private_start/end=313/313 exec=289 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X75:"xpc10:75" 1096 :  major_start_pcl=289   edge_private_start/end=312/312 exec=289 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X75:"xpc10:75" 1095 :  major_start_pcl=289   edge_private_start/end=311/311 exec=289 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X75:"xpc10:75" 1094 :  major_start_pcl=289   edge_private_start/end=310/310 exec=289 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X75:"xpc10:75" 1093 :  major_start_pcl=289   edge_private_start/end=309/309 exec=289 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X75:"xpc10:75" 1092 :  major_start_pcl=289   edge_private_start/end=308/308 exec=289 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X75:"xpc10:75" 1091 :  major_start_pcl=289   edge_private_start/end=307/307 exec=289 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X75:"xpc10:75" 1090 :  major_start_pcl=289   edge_private_start/end=306/306 exec=289 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X75:"xpc10:75" 1089 :  major_start_pcl=289   edge_private_start/end=305/305 exec=289 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X75:"xpc10:75" 1088 :  major_start_pcl=289   edge_private_start/end=304/304 exec=289 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X75:"xpc10:75" 1087 :  major_start_pcl=289   edge_private_start/end=303/303 exec=289 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X75:"xpc10:75" 1086 :  major_start_pcl=289   edge_private_start/end=302/302 exec=289 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X75:"xpc10:75" 1085 :  major_start_pcl=289   edge_private_start/end=301/301 exec=289 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X75:"xpc10:75" 1084 :  major_start_pcl=289   edge_private_start/end=300/300 exec=289 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X75:"xpc10:75" 1083 :  major_start_pcl=289   edge_private_start/end=299/299 exec=289 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X75:"xpc10:75" 1082 :  major_start_pcl=289   edge_private_start/end=298/298 exec=289 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X75:"xpc10:75" 1081 :  major_start_pcl=289   edge_private_start/end=297/297 exec=289 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X75:"xpc10:75" 1080 :  major_start_pcl=289   edge_private_start/end=296/296 exec=289 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X75:"xpc10:75" 1079 :  major_start_pcl=289   edge_private_start/end=295/295 exec=289 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X75:"xpc10:75" 1078 :  major_start_pcl=289   edge_private_start/end=294/294 exec=289 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X75:"xpc10:75" 1077 :  major_start_pcl=289   edge_private_start/end=293/293 exec=289 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X75:"xpc10:75" 1076 :  major_start_pcl=289   edge_private_start/end=292/292 exec=289 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X75:"xpc10:75" 1075 :  major_start_pcl=289   edge_private_start/end=291/291 exec=289 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X75:"xpc10:75" 1074 :  major_start_pcl=289   edge_private_start/end=290/290 exec=289 (dend=1)
//Simple greedy schedule for res2: Thread=xpc10 state=X75:"xpc10:75"
//res2: Thread=xpc10 state=X75:"xpc10:75"
//*-------+------+---------+-------------------------------------------------------------------------------------------------------------------------------------------------*
//| pc    | eno  | Phaser  | Work                                                                                                                                            |
//*-------+------+---------+-------------------------------------------------------------------------------------------------------------------------------------------------*
//| 289   | -    | R0 CTRL |                                                                                                                                                 |
//| 289   | 1074 | R0 DATA |                                                                                                                                                 |
//| 289+E | 1074 | W0 DATA | @_SINT/CC/MAPR10NoCE3_ARA0 te=te:289 write(TCin1.9_V_5, C(TCin1.9_V_0)) @_SINT/CC/MAPR12NoCE3_ARB0 te=te:289 write(TCin1.9_V_5, C(TCin1.9_V_2)) |
//| 290   | 1074 | W1 DATA |                                                                                                                                                 |
//| 289   | 1075 | R0 DATA |                                                                                                                                                 |
//| 289+E | 1075 | W0 DATA | @_SINT/CC/MAPR10NoCE3_ARA0 te=te:289 write(TCin1.9_V_5, C(TCin1.9_V_0)) @_SINT/CC/MAPR12NoCE2_ARB0 te=te:289 write(TCin1.9_V_5, C(TCin1.9_V_2)) |
//| 291   | 1075 | W1 DATA |                                                                                                                                                 |
//| 289   | 1076 | R0 DATA |                                                                                                                                                 |
//| 289+E | 1076 | W0 DATA | @_SINT/CC/MAPR10NoCE3_ARA0 te=te:289 write(TCin1.9_V_5, C(TCin1.9_V_0)) @_SINT/CC/MAPR12NoCE1_ARB0 te=te:289 write(TCin1.9_V_5, C(TCin1.9_V_2)) |
//| 292   | 1076 | W1 DATA |                                                                                                                                                 |
//| 289   | 1077 | R0 DATA |                                                                                                                                                 |
//| 289+E | 1077 | W0 DATA | @_SINT/CC/MAPR10NoCE3_ARA0 te=te:289 write(TCin1.9_V_5, C(TCin1.9_V_0)) @_SINT/CC/MAPR12NoCE0_ARB0 te=te:289 write(TCin1.9_V_5, C(TCin1.9_V_2)) |
//| 293   | 1077 | W1 DATA |                                                                                                                                                 |
//| 289   | 1078 | R0 DATA |                                                                                                                                                 |
//| 289+E | 1078 | W0 DATA | @_SINT/CC/MAPR10NoCE3_ARA0 te=te:289 write(TCin1.9_V_5, C(TCin1.9_V_0)) TCin1.9_V_0 te=te:289 scalarw(C(TCin1.9_V_6))                           |
//| 294   | 1078 | W1 DATA |                                                                                                                                                 |
//| 289   | 1079 | R0 DATA |                                                                                                                                                 |
//| 289+E | 1079 | W0 DATA | @_SINT/CC/MAPR10NoCE2_ARA0 te=te:289 write(TCin1.9_V_5, C(TCin1.9_V_0)) @_SINT/CC/MAPR12NoCE3_ARB0 te=te:289 write(TCin1.9_V_5, C(TCin1.9_V_2)) |
//| 295   | 1079 | W1 DATA |                                                                                                                                                 |
//| 289   | 1080 | R0 DATA |                                                                                                                                                 |
//| 289+E | 1080 | W0 DATA | @_SINT/CC/MAPR10NoCE2_ARA0 te=te:289 write(TCin1.9_V_5, C(TCin1.9_V_0)) @_SINT/CC/MAPR12NoCE2_ARB0 te=te:289 write(TCin1.9_V_5, C(TCin1.9_V_2)) |
//| 296   | 1080 | W1 DATA |                                                                                                                                                 |
//| 289   | 1081 | R0 DATA |                                                                                                                                                 |
//| 289+E | 1081 | W0 DATA | @_SINT/CC/MAPR10NoCE2_ARA0 te=te:289 write(TCin1.9_V_5, C(TCin1.9_V_0)) @_SINT/CC/MAPR12NoCE1_ARB0 te=te:289 write(TCin1.9_V_5, C(TCin1.9_V_2)) |
//| 297   | 1081 | W1 DATA |                                                                                                                                                 |
//| 289   | 1082 | R0 DATA |                                                                                                                                                 |
//| 289+E | 1082 | W0 DATA | @_SINT/CC/MAPR10NoCE2_ARA0 te=te:289 write(TCin1.9_V_5, C(TCin1.9_V_0)) @_SINT/CC/MAPR12NoCE0_ARB0 te=te:289 write(TCin1.9_V_5, C(TCin1.9_V_2)) |
//| 298   | 1082 | W1 DATA |                                                                                                                                                 |
//| 289   | 1083 | R0 DATA |                                                                                                                                                 |
//| 289+E | 1083 | W0 DATA | @_SINT/CC/MAPR10NoCE2_ARA0 te=te:289 write(TCin1.9_V_5, C(TCin1.9_V_0)) TCin1.9_V_0 te=te:289 scalarw(C(TCin1.9_V_6))                           |
//| 299   | 1083 | W1 DATA |                                                                                                                                                 |
//| 289   | 1084 | R0 DATA |                                                                                                                                                 |
//| 289+E | 1084 | W0 DATA | @_SINT/CC/MAPR10NoCE1_ARA0 te=te:289 write(TCin1.9_V_5, C(TCin1.9_V_0)) @_SINT/CC/MAPR12NoCE3_ARB0 te=te:289 write(TCin1.9_V_5, C(TCin1.9_V_2)) |
//| 300   | 1084 | W1 DATA |                                                                                                                                                 |
//| 289   | 1085 | R0 DATA |                                                                                                                                                 |
//| 289+E | 1085 | W0 DATA | @_SINT/CC/MAPR10NoCE1_ARA0 te=te:289 write(TCin1.9_V_5, C(TCin1.9_V_0)) @_SINT/CC/MAPR12NoCE2_ARB0 te=te:289 write(TCin1.9_V_5, C(TCin1.9_V_2)) |
//| 301   | 1085 | W1 DATA |                                                                                                                                                 |
//| 289   | 1086 | R0 DATA |                                                                                                                                                 |
//| 289+E | 1086 | W0 DATA | @_SINT/CC/MAPR10NoCE1_ARA0 te=te:289 write(TCin1.9_V_5, C(TCin1.9_V_0)) @_SINT/CC/MAPR12NoCE1_ARB0 te=te:289 write(TCin1.9_V_5, C(TCin1.9_V_2)) |
//| 302   | 1086 | W1 DATA |                                                                                                                                                 |
//| 289   | 1087 | R0 DATA |                                                                                                                                                 |
//| 289+E | 1087 | W0 DATA | @_SINT/CC/MAPR10NoCE1_ARA0 te=te:289 write(TCin1.9_V_5, C(TCin1.9_V_0)) @_SINT/CC/MAPR12NoCE0_ARB0 te=te:289 write(TCin1.9_V_5, C(TCin1.9_V_2)) |
//| 303   | 1087 | W1 DATA |                                                                                                                                                 |
//| 289   | 1088 | R0 DATA |                                                                                                                                                 |
//| 289+E | 1088 | W0 DATA | @_SINT/CC/MAPR10NoCE1_ARA0 te=te:289 write(TCin1.9_V_5, C(TCin1.9_V_0)) TCin1.9_V_0 te=te:289 scalarw(C(TCin1.9_V_6))                           |
//| 304   | 1088 | W1 DATA |                                                                                                                                                 |
//| 289   | 1089 | R0 DATA |                                                                                                                                                 |
//| 289+E | 1089 | W0 DATA | @_SINT/CC/MAPR10NoCE0_ARA0 te=te:289 write(TCin1.9_V_5, C(TCin1.9_V_0)) @_SINT/CC/MAPR12NoCE3_ARB0 te=te:289 write(TCin1.9_V_5, C(TCin1.9_V_2)) |
//| 305   | 1089 | W1 DATA |                                                                                                                                                 |
//| 289   | 1090 | R0 DATA |                                                                                                                                                 |
//| 289+E | 1090 | W0 DATA | @_SINT/CC/MAPR10NoCE0_ARA0 te=te:289 write(TCin1.9_V_5, C(TCin1.9_V_0)) @_SINT/CC/MAPR12NoCE2_ARB0 te=te:289 write(TCin1.9_V_5, C(TCin1.9_V_2)) |
//| 306   | 1090 | W1 DATA |                                                                                                                                                 |
//| 289   | 1091 | R0 DATA |                                                                                                                                                 |
//| 289+E | 1091 | W0 DATA | @_SINT/CC/MAPR10NoCE0_ARA0 te=te:289 write(TCin1.9_V_5, C(TCin1.9_V_0)) @_SINT/CC/MAPR12NoCE1_ARB0 te=te:289 write(TCin1.9_V_5, C(TCin1.9_V_2)) |
//| 307   | 1091 | W1 DATA |                                                                                                                                                 |
//| 289   | 1092 | R0 DATA |                                                                                                                                                 |
//| 289+E | 1092 | W0 DATA | @_SINT/CC/MAPR10NoCE0_ARA0 te=te:289 write(TCin1.9_V_5, C(TCin1.9_V_0)) @_SINT/CC/MAPR12NoCE0_ARB0 te=te:289 write(TCin1.9_V_5, C(TCin1.9_V_2)) |
//| 308   | 1092 | W1 DATA |                                                                                                                                                 |
//| 289   | 1093 | R0 DATA |                                                                                                                                                 |
//| 289+E | 1093 | W0 DATA | @_SINT/CC/MAPR10NoCE0_ARA0 te=te:289 write(TCin1.9_V_5, C(TCin1.9_V_0)) TCin1.9_V_0 te=te:289 scalarw(C(TCin1.9_V_6))                           |
//| 309   | 1093 | W1 DATA |                                                                                                                                                 |
//| 289   | 1094 | R0 DATA |                                                                                                                                                 |
//| 289+E | 1094 | W0 DATA | @_SINT/CC/MAPR12NoCE3_ARB0 te=te:289 write(TCin1.9_V_5, C(TCin1.9_V_2)) TCin1.9_V_0 te=te:289 scalarw(C(TCin1.9_V_6))                           |
//| 310   | 1094 | W1 DATA |                                                                                                                                                 |
//| 289   | 1095 | R0 DATA |                                                                                                                                                 |
//| 289+E | 1095 | W0 DATA | @_SINT/CC/MAPR12NoCE2_ARB0 te=te:289 write(TCin1.9_V_5, C(TCin1.9_V_2)) TCin1.9_V_0 te=te:289 scalarw(C(TCin1.9_V_6))                           |
//| 311   | 1095 | W1 DATA |                                                                                                                                                 |
//| 289   | 1096 | R0 DATA |                                                                                                                                                 |
//| 289+E | 1096 | W0 DATA | @_SINT/CC/MAPR12NoCE1_ARB0 te=te:289 write(TCin1.9_V_5, C(TCin1.9_V_2)) TCin1.9_V_0 te=te:289 scalarw(C(TCin1.9_V_6))                           |
//| 312   | 1096 | W1 DATA |                                                                                                                                                 |
//| 289   | 1097 | R0 DATA |                                                                                                                                                 |
//| 289+E | 1097 | W0 DATA | @_SINT/CC/MAPR12NoCE0_ARB0 te=te:289 write(TCin1.9_V_5, C(TCin1.9_V_2)) TCin1.9_V_0 te=te:289 scalarw(C(TCin1.9_V_6))                           |
//| 313   | 1097 | W1 DATA |                                                                                                                                                 |
//| 289   | 1098 | R0 DATA |                                                                                                                                                 |
//| 289+E | 1098 | W0 DATA | TCin1.9_V_0 te=te:289 scalarw(C(TCin1.9_V_6)) TCin1.9_V_2 te=te:289 scalarw(C(TCin1.9_V_7))                                                     |
//*-------+------+---------+-------------------------------------------------------------------------------------------------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X76:"xpc10:76" 1102 :  major_start_pcl=314   edge_private_start/end=-1/-1 exec=314 (dend=0)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X76:"xpc10:76" 1101 :  major_start_pcl=314   edge_private_start/end=317/317 exec=314 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X76:"xpc10:76" 1100 :  major_start_pcl=314   edge_private_start/end=316/316 exec=314 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X76:"xpc10:76" 1099 :  major_start_pcl=314   edge_private_start/end=315/315 exec=314 (dend=1)
//Simple greedy schedule for res2: Thread=xpc10 state=X76:"xpc10:76"
//res2: Thread=xpc10 state=X76:"xpc10:76"
//*-------+------+---------+-----------------------------------------------------------------------------------------------------------------------*
//| pc    | eno  | Phaser  | Work                                                                                                                  |
//*-------+------+---------+-----------------------------------------------------------------------------------------------------------------------*
//| 314   | -    | R0 CTRL |                                                                                                                       |
//| 314   | 1099 | R0 DATA |                                                                                                                       |
//| 314+E | 1099 | W0 DATA | @_SINT/CC/MAPR12NoCE2_ARB0 te=te:314 write(TCin1.9_V_5, C(TCin1.9_V_2)) TCin1.9_V_0 te=te:314 scalarw(C(TCin1.9_V_6)) |
//| 315   | 1099 | W1 DATA |                                                                                                                       |
//| 314   | 1100 | R0 DATA |                                                                                                                       |
//| 314+E | 1100 | W0 DATA | @_SINT/CC/MAPR12NoCE1_ARB0 te=te:314 write(TCin1.9_V_5, C(TCin1.9_V_2)) TCin1.9_V_0 te=te:314 scalarw(C(TCin1.9_V_6)) |
//| 316   | 1100 | W1 DATA |                                                                                                                       |
//| 314   | 1101 | R0 DATA |                                                                                                                       |
//| 314+E | 1101 | W0 DATA | @_SINT/CC/MAPR12NoCE0_ARB0 te=te:314 write(TCin1.9_V_5, C(TCin1.9_V_2)) TCin1.9_V_0 te=te:314 scalarw(C(TCin1.9_V_6)) |
//| 317   | 1101 | W1 DATA |                                                                                                                       |
//| 314   | 1102 | R0 DATA |                                                                                                                       |
//| 314+E | 1102 | W0 DATA | TCin1.9_V_0 te=te:314 scalarw(C(TCin1.9_V_6)) TCin1.9_V_2 te=te:314 scalarw(C(TCin1.9_V_7))                           |
//*-------+------+---------+-----------------------------------------------------------------------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X77:"xpc10:77" 1103 :  major_start_pcl=318   edge_private_start/end=-1/-1 exec=318 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X77:"xpc10:77"
//res2: Thread=xpc10 state=X77:"xpc10:77"
//*-------+------+---------+-----------------------------------------------*
//| pc    | eno  | Phaser  | Work                                          |
//*-------+------+---------+-----------------------------------------------*
//| 318   | -    | R0 CTRL |                                               |
//| 318   | 1103 | R0 DATA |                                               |
//| 318+E | 1103 | W0 DATA | TCin1.9_V_2 te=te:318 scalarw(C(TCin1.9_V_7)) |
//*-------+------+---------+-----------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X78:"xpc10:78" 1104 :  major_start_pcl=319   edge_private_start/end=-1/-1 exec=319 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X78:"xpc10:78"
//res2: Thread=xpc10 state=X78:"xpc10:78"
//*-------+------+---------+---------------------------------------*
//| pc    | eno  | Phaser  | Work                                  |
//*-------+------+---------+---------------------------------------*
//| 319   | -    | R0 CTRL |                                       |
//| 319   | 1104 | R0 DATA |                                       |
//| 319+E | 1104 | W0 DATA | fastspilldup26 te=te:319 scalarw(E17) |
//*-------+------+---------+---------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X79:"xpc10:79" 1105 :  major_start_pcl=320   edge_private_start/end=-1/-1 exec=320 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X79:"xpc10:79"
//res2: Thread=xpc10 state=X79:"xpc10:79"
//*-------+------+---------+----------------------------------------------------------------------------------------------------------------------*
//| pc    | eno  | Phaser  | Work                                                                                                                 |
//*-------+------+---------+----------------------------------------------------------------------------------------------------------------------*
//| 320   | -    | R0 CTRL |                                                                                                                      |
//| 320   | 1105 | R0 DATA |                                                                                                                      |
//| 320+E | 1105 | W0 DATA | TCin1.9_V_3 te=te:320 scalarw(C(fastspilldup26)) @_SINT/CC/SCALbx24_next_victim te=te:320 scalarw(C(fastspilldup26)) |
//*-------+------+---------+----------------------------------------------------------------------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X80:"xpc10:80" 1106 :  major_start_pcl=321   edge_private_start/end=-1/-1 exec=321 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X80:"xpc10:80"
//res2: Thread=xpc10 state=X80:"xpc10:80"
//*-------+------+---------+-----------------------------------------------------------------*
//| pc    | eno  | Phaser  | Work                                                            |
//*-------+------+---------+-----------------------------------------------------------------*
//| 321   | -    | R0 CTRL |                                                                 |
//| 321   | 1106 | R0 DATA |                                                                 |
//| 321+E | 1106 | W0 DATA | @_SINT/CC/SCALbx24_next_victim te=te:321 scalarw(TCin1.9_V_3%4) |
//*-------+------+---------+-----------------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X81:"xpc10:81" 1107 :  major_start_pcl=322   edge_private_start/end=-1/-1 exec=322 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X81:"xpc10:81"
//res2: Thread=xpc10 state=X81:"xpc10:81"
//*-------+------+---------+-------------------------------------------------------------------*
//| pc    | eno  | Phaser  | Work                                                              |
//*-------+------+---------+-------------------------------------------------------------------*
//| 322   | -    | R0 CTRL |                                                                   |
//| 322   | 1107 | R0 DATA |                                                                   |
//| 322+E | 1107 | W0 DATA | TCin1.9_V_4 te=te:322 scalarw(0) TCin1.9_V_5 te=te:322 scalarw(0) |
//*-------+------+---------+-------------------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X82:"xpc10:82" 1108 :  major_start_pcl=323   edge_private_start/end=-1/-1 exec=323 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X82:"xpc10:82"
//res2: Thread=xpc10 state=X82:"xpc10:82"
//*-------+------+---------+---------------------------------------*
//| pc    | eno  | Phaser  | Work                                  |
//*-------+------+---------+---------------------------------------*
//| 323   | -    | R0 CTRL |                                       |
//| 323   | 1108 | R0 DATA |                                       |
//| 323+E | 1108 | W0 DATA | fastspilldup26 te=te:323 scalarw(E17) |
//*-------+------+---------+---------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X83:"xpc10:83" 1111 :  major_start_pcl=324   edge_private_start/end=-1/-1 exec=324 (dend=0)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X83:"xpc10:83" 1110 :  major_start_pcl=324   edge_private_start/end=326/326 exec=324 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X83:"xpc10:83" 1109 :  major_start_pcl=324   edge_private_start/end=325/325 exec=324 (dend=1)
//Simple greedy schedule for res2: Thread=xpc10 state=X83:"xpc10:83"
//res2: Thread=xpc10 state=X83:"xpc10:83"
//*-------+------+---------+-----------------------------------------------------------------------------------------------------------------------*
//| pc    | eno  | Phaser  | Work                                                                                                                  |
//*-------+------+---------+-----------------------------------------------------------------------------------------------------------------------*
//| 324   | -    | R0 CTRL |                                                                                                                       |
//| 324   | 1109 | R0 DATA |                                                                                                                       |
//| 324+E | 1109 | W0 DATA | @_SINT/CC/MAPR12NoCE1_ARB0 te=te:324 write(TCin1.9_V_5, C(TCin1.9_V_2)) TCin1.9_V_0 te=te:324 scalarw(C(TCin1.9_V_6)) |
//| 325   | 1109 | W1 DATA |                                                                                                                       |
//| 324   | 1110 | R0 DATA |                                                                                                                       |
//| 324+E | 1110 | W0 DATA | @_SINT/CC/MAPR12NoCE0_ARB0 te=te:324 write(TCin1.9_V_5, C(TCin1.9_V_2)) TCin1.9_V_0 te=te:324 scalarw(C(TCin1.9_V_6)) |
//| 326   | 1110 | W1 DATA |                                                                                                                       |
//| 324   | 1111 | R0 DATA |                                                                                                                       |
//| 324+E | 1111 | W0 DATA | TCin1.9_V_0 te=te:324 scalarw(C(TCin1.9_V_6)) TCin1.9_V_2 te=te:324 scalarw(C(TCin1.9_V_7))                           |
//*-------+------+---------+-----------------------------------------------------------------------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X84:"xpc10:84" 1113 :  major_start_pcl=327   edge_private_start/end=-1/-1 exec=327 (dend=0)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X84:"xpc10:84" 1112 :  major_start_pcl=327   edge_private_start/end=328/328 exec=327 (dend=1)
//Simple greedy schedule for res2: Thread=xpc10 state=X84:"xpc10:84"
//res2: Thread=xpc10 state=X84:"xpc10:84"
//*-------+------+---------+-----------------------------------------------------------------------------------------------------------------------*
//| pc    | eno  | Phaser  | Work                                                                                                                  |
//*-------+------+---------+-----------------------------------------------------------------------------------------------------------------------*
//| 327   | -    | R0 CTRL |                                                                                                                       |
//| 327   | 1112 | R0 DATA |                                                                                                                       |
//| 327+E | 1112 | W0 DATA | @_SINT/CC/MAPR12NoCE0_ARB0 te=te:327 write(TCin1.9_V_5, C(TCin1.9_V_2)) TCin1.9_V_0 te=te:327 scalarw(C(TCin1.9_V_6)) |
//| 328   | 1112 | W1 DATA |                                                                                                                       |
//| 327   | 1113 | R0 DATA |                                                                                                                       |
//| 327+E | 1113 | W0 DATA | TCin1.9_V_0 te=te:327 scalarw(C(TCin1.9_V_6)) TCin1.9_V_2 te=te:327 scalarw(C(TCin1.9_V_7))                           |
//*-------+------+---------+-----------------------------------------------------------------------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X85:"xpc10:85" 1114 :  major_start_pcl=329   edge_private_start/end=-1/-1 exec=329 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X85:"xpc10:85"
//res2: Thread=xpc10 state=X85:"xpc10:85"
//*-------+------+---------+---------------------------------------------------------------------------------------------*
//| pc    | eno  | Phaser  | Work                                                                                        |
//*-------+------+---------+---------------------------------------------------------------------------------------------*
//| 329   | -    | R0 CTRL |                                                                                             |
//| 329   | 1114 | R0 DATA |                                                                                             |
//| 329+E | 1114 | W0 DATA | TCin1.9_V_0 te=te:329 scalarw(C(TCin1.9_V_6)) TCin1.9_V_2 te=te:329 scalarw(C(TCin1.9_V_7)) |
//*-------+------+---------+---------------------------------------------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X86:"xpc10:86" 1118 :  major_start_pcl=330   edge_private_start/end=-1/-1 exec=330 (dend=0)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X86:"xpc10:86" 1117 :  major_start_pcl=330   edge_private_start/end=333/333 exec=330 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X86:"xpc10:86" 1116 :  major_start_pcl=330   edge_private_start/end=332/332 exec=330 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X86:"xpc10:86" 1115 :  major_start_pcl=330   edge_private_start/end=331/331 exec=330 (dend=1)
//Simple greedy schedule for res2: Thread=xpc10 state=X86:"xpc10:86"
//res2: Thread=xpc10 state=X86:"xpc10:86"
//*-------+------+---------+--------------------------------------------------------------------------------------------------------------*
//| pc    | eno  | Phaser  | Work                                                                                                         |
//*-------+------+---------+--------------------------------------------------------------------------------------------------------------*
//| 330   | -    | R0 CTRL |                                                                                                              |
//| 330   | 1115 | R0 DATA |                                                                                                              |
//| 330+E | 1115 | W0 DATA | @_SINT/CC/MAPR12NoCE2_ARB0 te=te:330 write(TCin1.9_V_5, C(TCin1.9_V_2)) TCi1._SPILL_256 te=te:330 scalarw(0) |
//| 331   | 1115 | W1 DATA |                                                                                                              |
//| 330   | 1116 | R0 DATA |                                                                                                              |
//| 330+E | 1116 | W0 DATA | @_SINT/CC/MAPR12NoCE1_ARB0 te=te:330 write(TCin1.9_V_5, C(TCin1.9_V_2)) TCi1._SPILL_256 te=te:330 scalarw(0) |
//| 332   | 1116 | W1 DATA |                                                                                                              |
//| 330   | 1117 | R0 DATA |                                                                                                              |
//| 330+E | 1117 | W0 DATA | @_SINT/CC/MAPR12NoCE0_ARB0 te=te:330 write(TCin1.9_V_5, C(TCin1.9_V_2)) TCi1._SPILL_256 te=te:330 scalarw(0) |
//| 333   | 1117 | W1 DATA |                                                                                                              |
//| 330   | 1118 | R0 DATA |                                                                                                              |
//| 330+E | 1118 | W0 DATA | TTMT4Main_V_7 te=te:330 scalarw(S32'0I) TCi1._SPILL_256 te=te:330 scalarw(0)                                 |
//*-------+------+---------+--------------------------------------------------------------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X87:"xpc10:87" 1120 :  major_start_pcl=334   edge_private_start/end=-1/-1 exec=334 (dend=0)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X87:"xpc10:87" 1119 :  major_start_pcl=334   edge_private_start/end=-1/-1 exec=334 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X87:"xpc10:87"
//res2: Thread=xpc10 state=X87:"xpc10:87"
//*-------+------+---------+------------------------------------------------------------------------------------------------------*
//| pc    | eno  | Phaser  | Work                                                                                                 |
//*-------+------+---------+------------------------------------------------------------------------------------------------------*
//| 334   | -    | R0 CTRL |                                                                                                      |
//| 334   | 1119 | R0 DATA |                                                                                                      |
//| 334+E | 1119 | W0 DATA | TTMT4Main_V_3 te=te:334 scalarw(1+TTMT4Main_V_3) TTMT4Main_V_7 te=te:334 scalarw(C(TCi1._SPILL_256)) |
//| 334   | 1120 | R0 DATA |                                                                                                      |
//| 334+E | 1120 | W0 DATA | TTMT4Main_V_2 te=te:334 scalarw(1+TTMT4Main_V_2) TTMT4Main_V_7 te=te:334 scalarw(C(TCi1._SPILL_256)) |
//*-------+------+---------+------------------------------------------------------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X88:"xpc10:88" 1123 :  major_start_pcl=335   edge_private_start/end=-1/-1 exec=335 (dend=0)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X88:"xpc10:88" 1122 :  major_start_pcl=335   edge_private_start/end=337/337 exec=335 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X88:"xpc10:88" 1121 :  major_start_pcl=335   edge_private_start/end=336/336 exec=335 (dend=1)
//Simple greedy schedule for res2: Thread=xpc10 state=X88:"xpc10:88"
//res2: Thread=xpc10 state=X88:"xpc10:88"
//*-------+------+---------+--------------------------------------------------------------------------------------------------------------*
//| pc    | eno  | Phaser  | Work                                                                                                         |
//*-------+------+---------+--------------------------------------------------------------------------------------------------------------*
//| 335   | -    | R0 CTRL |                                                                                                              |
//| 335   | 1121 | R0 DATA |                                                                                                              |
//| 335+E | 1121 | W0 DATA | @_SINT/CC/MAPR12NoCE1_ARB0 te=te:335 write(TCin1.9_V_5, C(TCin1.9_V_2)) TCi1._SPILL_256 te=te:335 scalarw(0) |
//| 336   | 1121 | W1 DATA |                                                                                                              |
//| 335   | 1122 | R0 DATA |                                                                                                              |
//| 335+E | 1122 | W0 DATA | @_SINT/CC/MAPR12NoCE0_ARB0 te=te:335 write(TCin1.9_V_5, C(TCin1.9_V_2)) TCi1._SPILL_256 te=te:335 scalarw(0) |
//| 337   | 1122 | W1 DATA |                                                                                                              |
//| 335   | 1123 | R0 DATA |                                                                                                              |
//| 335+E | 1123 | W0 DATA | TTMT4Main_V_7 te=te:335 scalarw(S32'0I) TCi1._SPILL_256 te=te:335 scalarw(0)                                 |
//*-------+------+---------+--------------------------------------------------------------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X89:"xpc10:89" 1125 :  major_start_pcl=338   edge_private_start/end=-1/-1 exec=338 (dend=0)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X89:"xpc10:89" 1124 :  major_start_pcl=338   edge_private_start/end=339/339 exec=338 (dend=1)
//Simple greedy schedule for res2: Thread=xpc10 state=X89:"xpc10:89"
//res2: Thread=xpc10 state=X89:"xpc10:89"
//*-------+------+---------+--------------------------------------------------------------------------------------------------------------*
//| pc    | eno  | Phaser  | Work                                                                                                         |
//*-------+------+---------+--------------------------------------------------------------------------------------------------------------*
//| 338   | -    | R0 CTRL |                                                                                                              |
//| 338   | 1124 | R0 DATA |                                                                                                              |
//| 338+E | 1124 | W0 DATA | @_SINT/CC/MAPR12NoCE0_ARB0 te=te:338 write(TCin1.9_V_5, C(TCin1.9_V_2)) TCi1._SPILL_256 te=te:338 scalarw(0) |
//| 339   | 1124 | W1 DATA |                                                                                                              |
//| 338   | 1125 | R0 DATA |                                                                                                              |
//| 338+E | 1125 | W0 DATA | TTMT4Main_V_7 te=te:338 scalarw(S32'0I) TCi1._SPILL_256 te=te:338 scalarw(0)                                 |
//*-------+------+---------+--------------------------------------------------------------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X90:"xpc10:90" 1126 :  major_start_pcl=340   edge_private_start/end=-1/-1 exec=340 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X90:"xpc10:90"
//res2: Thread=xpc10 state=X90:"xpc10:90"
//*-------+------+---------+------------------------------------------------------------------------------*
//| pc    | eno  | Phaser  | Work                                                                         |
//*-------+------+---------+------------------------------------------------------------------------------*
//| 340   | -    | R0 CTRL |                                                                              |
//| 340   | 1126 | R0 DATA |                                                                              |
//| 340+E | 1126 | W0 DATA | TTMT4Main_V_7 te=te:340 scalarw(S32'0I) TCi1._SPILL_256 te=te:340 scalarw(0) |
//*-------+------+---------+------------------------------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X91:"xpc10:91" 1127 :  major_start_pcl=341   edge_private_start/end=-1/-1 exec=341 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X91:"xpc10:91"
//res2: Thread=xpc10 state=X91:"xpc10:91"
//*-------+------+---------+-------------------------------------*
//| pc    | eno  | Phaser  | Work                                |
//*-------+------+---------+-------------------------------------*
//| 341   | -    | R0 CTRL |                                     |
//| 341   | 1127 | R0 DATA |                                     |
//| 341+E | 1127 | W0 DATA | TCha6.10_V_0 te=te:341 scalarw(E18) |
//*-------+------+---------+-------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X92:"xpc10:92" 1129 :  major_start_pcl=342   edge_private_start/end=343/406 exec=406 (dend=64)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X92:"xpc10:92" 1128 :  major_start_pcl=342   edge_private_start/end=-1/-1 exec=342 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X92:"xpc10:92"
//res2: Thread=xpc10 state=X92:"xpc10:92"
//*---------+------+----------+----------------------------------------------------------*
//| pc      | eno  | Phaser   | Work                                                     |
//*---------+------+----------+----------------------------------------------------------*
//| 342     | -    | R0 CTRL  |                                                          |
//| 342     | 1128 | R0 DATA  |                                                          |
//| 342+E   | 1128 | W0 DATA  | TCha6.10_V_0 te=te:342 scalarw(-TCha6.10_V_0)            |
//| 342+S   | 1129 | R0 DATA  | isMODULUS10 te=te:342 *fixed-func-ALU*(TCha6.10_V_0, E7) |
//| 343     | 1129 | R1 DATA  |                                                          |
//| 344     | 1129 | R2 DATA  |                                                          |
//| 345     | 1129 | R3 DATA  |                                                          |
//| 346     | 1129 | R4 DATA  |                                                          |
//| 347     | 1129 | R5 DATA  |                                                          |
//| 348     | 1129 | R6 DATA  |                                                          |
//| 349     | 1129 | R7 DATA  |                                                          |
//| 350     | 1129 | R8 DATA  |                                                          |
//| 351     | 1129 | R9 DATA  |                                                          |
//| 352     | 1129 | R10 DATA |                                                          |
//| 353     | 1129 | R11 DATA |                                                          |
//| 354     | 1129 | R12 DATA |                                                          |
//| 355     | 1129 | R13 DATA |                                                          |
//| 356     | 1129 | R14 DATA |                                                          |
//| 357     | 1129 | R15 DATA |                                                          |
//| 358     | 1129 | R16 DATA |                                                          |
//| 359     | 1129 | R17 DATA |                                                          |
//| 360     | 1129 | R18 DATA |                                                          |
//| 361     | 1129 | R19 DATA |                                                          |
//| 362     | 1129 | R20 DATA |                                                          |
//| 363     | 1129 | R21 DATA |                                                          |
//| 364     | 1129 | R22 DATA |                                                          |
//| 365     | 1129 | R23 DATA |                                                          |
//| 366     | 1129 | R24 DATA |                                                          |
//| 367     | 1129 | R25 DATA |                                                          |
//| 368     | 1129 | R26 DATA |                                                          |
//| 369     | 1129 | R27 DATA |                                                          |
//| 370     | 1129 | R28 DATA |                                                          |
//| 371     | 1129 | R29 DATA |                                                          |
//| 372     | 1129 | R30 DATA |                                                          |
//| 373     | 1129 | R31 DATA |                                                          |
//| 374     | 1129 | R32 DATA |                                                          |
//| 375     | 1129 | R33 DATA |                                                          |
//| 376     | 1129 | R34 DATA |                                                          |
//| 377     | 1129 | R35 DATA |                                                          |
//| 378     | 1129 | R36 DATA |                                                          |
//| 379     | 1129 | R37 DATA |                                                          |
//| 380     | 1129 | R38 DATA |                                                          |
//| 381     | 1129 | R39 DATA |                                                          |
//| 382     | 1129 | R40 DATA |                                                          |
//| 383     | 1129 | R41 DATA |                                                          |
//| 384     | 1129 | R42 DATA |                                                          |
//| 385     | 1129 | R43 DATA |                                                          |
//| 386     | 1129 | R44 DATA |                                                          |
//| 387     | 1129 | R45 DATA |                                                          |
//| 388     | 1129 | R46 DATA |                                                          |
//| 389     | 1129 | R47 DATA |                                                          |
//| 390     | 1129 | R48 DATA |                                                          |
//| 391     | 1129 | R49 DATA |                                                          |
//| 392     | 1129 | R50 DATA |                                                          |
//| 393     | 1129 | R51 DATA |                                                          |
//| 394     | 1129 | R52 DATA |                                                          |
//| 395     | 1129 | R53 DATA |                                                          |
//| 396     | 1129 | R54 DATA |                                                          |
//| 397     | 1129 | R55 DATA |                                                          |
//| 398     | 1129 | R56 DATA |                                                          |
//| 399     | 1129 | R57 DATA |                                                          |
//| 400     | 1129 | R58 DATA |                                                          |
//| 401     | 1129 | R59 DATA |                                                          |
//| 402     | 1129 | R60 DATA |                                                          |
//| 403     | 1129 | R61 DATA |                                                          |
//| 404     | 1129 | R62 DATA |                                                          |
//| 405     | 1129 | R63 DATA |                                                          |
//| 406+S   | 1129 | R64 DATA |                                                          |
//| 406+E+S | 1129 | W0 DATA  | TCin1.9_V_5 te=te:406 scalarw(E19)                       |
//*---------+------+----------+----------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X93:"xpc10:93" 1130 :  major_start_pcl=407   edge_private_start/end=408/471 exec=471 (dend=64)
//Simple greedy schedule for res2: Thread=xpc10 state=X93:"xpc10:93"
//res2: Thread=xpc10 state=X93:"xpc10:93"
//*---------+------+----------+----------------------------------------------------------*
//| pc      | eno  | Phaser   | Work                                                     |
//*---------+------+----------+----------------------------------------------------------*
//| 407     | -    | R0 CTRL  |                                                          |
//| 407+S   | 1130 | R0 DATA  | isMODULUS10 te=te:407 *fixed-func-ALU*(TCha6.10_V_0, E7) |
//| 408     | 1130 | R1 DATA  |                                                          |
//| 409     | 1130 | R2 DATA  |                                                          |
//| 410     | 1130 | R3 DATA  |                                                          |
//| 411     | 1130 | R4 DATA  |                                                          |
//| 412     | 1130 | R5 DATA  |                                                          |
//| 413     | 1130 | R6 DATA  |                                                          |
//| 414     | 1130 | R7 DATA  |                                                          |
//| 415     | 1130 | R8 DATA  |                                                          |
//| 416     | 1130 | R9 DATA  |                                                          |
//| 417     | 1130 | R10 DATA |                                                          |
//| 418     | 1130 | R11 DATA |                                                          |
//| 419     | 1130 | R12 DATA |                                                          |
//| 420     | 1130 | R13 DATA |                                                          |
//| 421     | 1130 | R14 DATA |                                                          |
//| 422     | 1130 | R15 DATA |                                                          |
//| 423     | 1130 | R16 DATA |                                                          |
//| 424     | 1130 | R17 DATA |                                                          |
//| 425     | 1130 | R18 DATA |                                                          |
//| 426     | 1130 | R19 DATA |                                                          |
//| 427     | 1130 | R20 DATA |                                                          |
//| 428     | 1130 | R21 DATA |                                                          |
//| 429     | 1130 | R22 DATA |                                                          |
//| 430     | 1130 | R23 DATA |                                                          |
//| 431     | 1130 | R24 DATA |                                                          |
//| 432     | 1130 | R25 DATA |                                                          |
//| 433     | 1130 | R26 DATA |                                                          |
//| 434     | 1130 | R27 DATA |                                                          |
//| 435     | 1130 | R28 DATA |                                                          |
//| 436     | 1130 | R29 DATA |                                                          |
//| 437     | 1130 | R30 DATA |                                                          |
//| 438     | 1130 | R31 DATA |                                                          |
//| 439     | 1130 | R32 DATA |                                                          |
//| 440     | 1130 | R33 DATA |                                                          |
//| 441     | 1130 | R34 DATA |                                                          |
//| 442     | 1130 | R35 DATA |                                                          |
//| 443     | 1130 | R36 DATA |                                                          |
//| 444     | 1130 | R37 DATA |                                                          |
//| 445     | 1130 | R38 DATA |                                                          |
//| 446     | 1130 | R39 DATA |                                                          |
//| 447     | 1130 | R40 DATA |                                                          |
//| 448     | 1130 | R41 DATA |                                                          |
//| 449     | 1130 | R42 DATA |                                                          |
//| 450     | 1130 | R43 DATA |                                                          |
//| 451     | 1130 | R44 DATA |                                                          |
//| 452     | 1130 | R45 DATA |                                                          |
//| 453     | 1130 | R46 DATA |                                                          |
//| 454     | 1130 | R47 DATA |                                                          |
//| 455     | 1130 | R48 DATA |                                                          |
//| 456     | 1130 | R49 DATA |                                                          |
//| 457     | 1130 | R50 DATA |                                                          |
//| 458     | 1130 | R51 DATA |                                                          |
//| 459     | 1130 | R52 DATA |                                                          |
//| 460     | 1130 | R53 DATA |                                                          |
//| 461     | 1130 | R54 DATA |                                                          |
//| 462     | 1130 | R55 DATA |                                                          |
//| 463     | 1130 | R56 DATA |                                                          |
//| 464     | 1130 | R57 DATA |                                                          |
//| 465     | 1130 | R58 DATA |                                                          |
//| 466     | 1130 | R59 DATA |                                                          |
//| 467     | 1130 | R60 DATA |                                                          |
//| 468     | 1130 | R61 DATA |                                                          |
//| 469     | 1130 | R62 DATA |                                                          |
//| 470     | 1130 | R63 DATA |                                                          |
//| 471+S   | 1130 | R64 DATA |                                                          |
//| 471+E+S | 1130 | W0 DATA  | TCin1.9_V_5 te=te:471 scalarw(E19)                       |
//*---------+------+----------+----------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X94:"xpc10:94" 1161 :  major_start_pcl=472   edge_private_start/end=-1/-1 exec=473 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X94:"xpc10:94" 1160 :  major_start_pcl=472   edge_private_start/end=-1/-1 exec=473 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X94:"xpc10:94" 1159 :  major_start_pcl=472   edge_private_start/end=501/501 exec=473 (dend=2)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X94:"xpc10:94" 1158 :  major_start_pcl=472   edge_private_start/end=500/500 exec=473 (dend=2)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X94:"xpc10:94" 1157 :  major_start_pcl=472   edge_private_start/end=499/499 exec=473 (dend=2)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X94:"xpc10:94" 1156 :  major_start_pcl=472   edge_private_start/end=498/498 exec=473 (dend=2)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X94:"xpc10:94" 1155 :  major_start_pcl=472   edge_private_start/end=-1/-1 exec=473 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X94:"xpc10:94" 1154 :  major_start_pcl=472   edge_private_start/end=497/497 exec=473 (dend=2)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X94:"xpc10:94" 1153 :  major_start_pcl=472   edge_private_start/end=496/496 exec=473 (dend=2)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X94:"xpc10:94" 1152 :  major_start_pcl=472   edge_private_start/end=495/495 exec=473 (dend=2)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X94:"xpc10:94" 1151 :  major_start_pcl=472   edge_private_start/end=494/494 exec=473 (dend=2)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X94:"xpc10:94" 1150 :  major_start_pcl=472   edge_private_start/end=493/493 exec=473 (dend=2)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X94:"xpc10:94" 1149 :  major_start_pcl=472   edge_private_start/end=492/492 exec=473 (dend=2)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X94:"xpc10:94" 1148 :  major_start_pcl=472   edge_private_start/end=491/491 exec=473 (dend=2)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X94:"xpc10:94" 1147 :  major_start_pcl=472   edge_private_start/end=490/490 exec=473 (dend=2)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X94:"xpc10:94" 1146 :  major_start_pcl=472   edge_private_start/end=489/489 exec=473 (dend=2)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X94:"xpc10:94" 1145 :  major_start_pcl=472   edge_private_start/end=488/488 exec=473 (dend=2)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X94:"xpc10:94" 1144 :  major_start_pcl=472   edge_private_start/end=487/487 exec=473 (dend=2)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X94:"xpc10:94" 1143 :  major_start_pcl=472   edge_private_start/end=486/486 exec=473 (dend=2)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X94:"xpc10:94" 1142 :  major_start_pcl=472   edge_private_start/end=485/485 exec=473 (dend=2)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X94:"xpc10:94" 1141 :  major_start_pcl=472   edge_private_start/end=484/484 exec=473 (dend=2)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X94:"xpc10:94" 1140 :  major_start_pcl=472   edge_private_start/end=483/483 exec=473 (dend=2)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X94:"xpc10:94" 1139 :  major_start_pcl=472   edge_private_start/end=482/482 exec=473 (dend=2)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X94:"xpc10:94" 1138 :  major_start_pcl=472   edge_private_start/end=481/481 exec=473 (dend=2)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X94:"xpc10:94" 1137 :  major_start_pcl=472   edge_private_start/end=480/480 exec=473 (dend=2)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X94:"xpc10:94" 1136 :  major_start_pcl=472   edge_private_start/end=479/479 exec=473 (dend=2)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X94:"xpc10:94" 1135 :  major_start_pcl=472   edge_private_start/end=478/478 exec=473 (dend=2)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X94:"xpc10:94" 1134 :  major_start_pcl=472   edge_private_start/end=477/477 exec=473 (dend=2)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X94:"xpc10:94" 1133 :  major_start_pcl=472   edge_private_start/end=476/476 exec=473 (dend=2)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X94:"xpc10:94" 1132 :  major_start_pcl=472   edge_private_start/end=475/475 exec=473 (dend=2)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X94:"xpc10:94" 1131 :  major_start_pcl=472   edge_private_start/end=474/474 exec=473 (dend=2)
//Simple greedy schedule for res2: Thread=xpc10 state=X94:"xpc10:94"
//res2: Thread=xpc10 state=X94:"xpc10:94"
//*-------+------+---------+----------------------------------------------------------------------------------------------------------------------------------------------------*
//| pc    | eno  | Phaser  | Work                                                                                                                                               |
//*-------+------+---------+----------------------------------------------------------------------------------------------------------------------------------------------------*
//| 472   | -    | R0 CTRL | @_SINT/CC/MAPR10NoCE3_ARA0 te=te:472 read(TCin1.9_V_5) @_SINT/CC/MAPR10NoCE2_ARA0 te=te:472 read(TCin1.9_V_5) @_SINT/CC/MAPR10NoCE1_ARA0 te=te:47\ |
//|       |      |         | 2 read(TCin1.9_V_5) @_SINT/CC/MAPR10NoCE0_ARA0 te=te:472 read(TCin1.9_V_5)                                                                         |
//| 473   | -    | R1 CTRL |                                                                                                                                                    |
//| 472   | 1131 | R0 DATA |                                                                                                                                                    |
//| 473   | 1131 | R1 DATA |                                                                                                                                                    |
//| 473+E | 1131 | W0 DATA | @_SINT/CC/MAPR10NoCE3_ARA0 te=te:473 write(TCin1.9_V_5, C(TCin1.9_V_0))  PLI:Eviction %u needed                                                    |
//| 474   | 1131 | W1 DATA |                                                                                                                                                    |
//| 472   | 1132 | R0 DATA |                                                                                                                                                    |
//| 473   | 1132 | R1 DATA |                                                                                                                                                    |
//| 473+E | 1132 | W0 DATA | @_SINT/CC/MAPR10NoCE3_ARA0 te=te:473 write(TCin1.9_V_5, C(TCin1.9_V_0)) @_SINT/CC/MAPR12NoCE3_ARB0 te=te:473 write(TCin1.9_V_5, C(TCin1.9_V_2))    |
//| 475   | 1132 | W1 DATA |                                                                                                                                                    |
//| 472   | 1133 | R0 DATA |                                                                                                                                                    |
//| 473   | 1133 | R1 DATA |                                                                                                                                                    |
//| 473+E | 1133 | W0 DATA | @_SINT/CC/MAPR10NoCE3_ARA0 te=te:473 write(TCin1.9_V_5, C(TCin1.9_V_0)) @_SINT/CC/MAPR12NoCE2_ARB0 te=te:473 write(TCin1.9_V_5, C(TCin1.9_V_2))    |
//| 476   | 1133 | W1 DATA |                                                                                                                                                    |
//| 472   | 1134 | R0 DATA |                                                                                                                                                    |
//| 473   | 1134 | R1 DATA |                                                                                                                                                    |
//| 473+E | 1134 | W0 DATA | @_SINT/CC/MAPR10NoCE3_ARA0 te=te:473 write(TCin1.9_V_5, C(TCin1.9_V_0)) @_SINT/CC/MAPR12NoCE1_ARB0 te=te:473 write(TCin1.9_V_5, C(TCin1.9_V_2))    |
//| 477   | 1134 | W1 DATA |                                                                                                                                                    |
//| 472   | 1135 | R0 DATA |                                                                                                                                                    |
//| 473   | 1135 | R1 DATA |                                                                                                                                                    |
//| 473+E | 1135 | W0 DATA | @_SINT/CC/MAPR10NoCE3_ARA0 te=te:473 write(TCin1.9_V_5, C(TCin1.9_V_0)) @_SINT/CC/MAPR12NoCE0_ARB0 te=te:473 write(TCin1.9_V_5, C(TCin1.9_V_2))    |
//| 478   | 1135 | W1 DATA |                                                                                                                                                    |
//| 472   | 1136 | R0 DATA |                                                                                                                                                    |
//| 473   | 1136 | R1 DATA |                                                                                                                                                    |
//| 473+E | 1136 | W0 DATA | @_SINT/CC/MAPR10NoCE3_ARA0 te=te:473 write(TCin1.9_V_5, C(TCin1.9_V_0)) TCi1._SPILL_256 te=te:473 scalarw(0)                                       |
//| 479   | 1136 | W1 DATA |                                                                                                                                                    |
//| 472   | 1137 | R0 DATA |                                                                                                                                                    |
//| 473   | 1137 | R1 DATA |                                                                                                                                                    |
//| 473+E | 1137 | W0 DATA | @_SINT/CC/MAPR10NoCE2_ARA0 te=te:473 write(TCin1.9_V_5, C(TCin1.9_V_0))  PLI:Eviction %u needed                                                    |
//| 480   | 1137 | W1 DATA |                                                                                                                                                    |
//| 472   | 1138 | R0 DATA |                                                                                                                                                    |
//| 473   | 1138 | R1 DATA |                                                                                                                                                    |
//| 473+E | 1138 | W0 DATA | @_SINT/CC/MAPR10NoCE2_ARA0 te=te:473 write(TCin1.9_V_5, C(TCin1.9_V_0)) @_SINT/CC/MAPR12NoCE3_ARB0 te=te:473 write(TCin1.9_V_5, C(TCin1.9_V_2))    |
//| 481   | 1138 | W1 DATA |                                                                                                                                                    |
//| 472   | 1139 | R0 DATA |                                                                                                                                                    |
//| 473   | 1139 | R1 DATA |                                                                                                                                                    |
//| 473+E | 1139 | W0 DATA | @_SINT/CC/MAPR10NoCE2_ARA0 te=te:473 write(TCin1.9_V_5, C(TCin1.9_V_0)) @_SINT/CC/MAPR12NoCE2_ARB0 te=te:473 write(TCin1.9_V_5, C(TCin1.9_V_2))    |
//| 482   | 1139 | W1 DATA |                                                                                                                                                    |
//| 472   | 1140 | R0 DATA |                                                                                                                                                    |
//| 473   | 1140 | R1 DATA |                                                                                                                                                    |
//| 473+E | 1140 | W0 DATA | @_SINT/CC/MAPR10NoCE2_ARA0 te=te:473 write(TCin1.9_V_5, C(TCin1.9_V_0)) @_SINT/CC/MAPR12NoCE1_ARB0 te=te:473 write(TCin1.9_V_5, C(TCin1.9_V_2))    |
//| 483   | 1140 | W1 DATA |                                                                                                                                                    |
//| 472   | 1141 | R0 DATA |                                                                                                                                                    |
//| 473   | 1141 | R1 DATA |                                                                                                                                                    |
//| 473+E | 1141 | W0 DATA | @_SINT/CC/MAPR10NoCE2_ARA0 te=te:473 write(TCin1.9_V_5, C(TCin1.9_V_0)) @_SINT/CC/MAPR12NoCE0_ARB0 te=te:473 write(TCin1.9_V_5, C(TCin1.9_V_2))    |
//| 484   | 1141 | W1 DATA |                                                                                                                                                    |
//| 472   | 1142 | R0 DATA |                                                                                                                                                    |
//| 473   | 1142 | R1 DATA |                                                                                                                                                    |
//| 473+E | 1142 | W0 DATA | @_SINT/CC/MAPR10NoCE2_ARA0 te=te:473 write(TCin1.9_V_5, C(TCin1.9_V_0)) TCi1._SPILL_256 te=te:473 scalarw(0)                                       |
//| 485   | 1142 | W1 DATA |                                                                                                                                                    |
//| 472   | 1143 | R0 DATA |                                                                                                                                                    |
//| 473   | 1143 | R1 DATA |                                                                                                                                                    |
//| 473+E | 1143 | W0 DATA | @_SINT/CC/MAPR10NoCE1_ARA0 te=te:473 write(TCin1.9_V_5, C(TCin1.9_V_0))  PLI:Eviction %u needed                                                    |
//| 486   | 1143 | W1 DATA |                                                                                                                                                    |
//| 472   | 1144 | R0 DATA |                                                                                                                                                    |
//| 473   | 1144 | R1 DATA |                                                                                                                                                    |
//| 473+E | 1144 | W0 DATA | @_SINT/CC/MAPR10NoCE1_ARA0 te=te:473 write(TCin1.9_V_5, C(TCin1.9_V_0)) @_SINT/CC/MAPR12NoCE3_ARB0 te=te:473 write(TCin1.9_V_5, C(TCin1.9_V_2))    |
//| 487   | 1144 | W1 DATA |                                                                                                                                                    |
//| 472   | 1145 | R0 DATA |                                                                                                                                                    |
//| 473   | 1145 | R1 DATA |                                                                                                                                                    |
//| 473+E | 1145 | W0 DATA | @_SINT/CC/MAPR10NoCE1_ARA0 te=te:473 write(TCin1.9_V_5, C(TCin1.9_V_0)) @_SINT/CC/MAPR12NoCE2_ARB0 te=te:473 write(TCin1.9_V_5, C(TCin1.9_V_2))    |
//| 488   | 1145 | W1 DATA |                                                                                                                                                    |
//| 472   | 1146 | R0 DATA |                                                                                                                                                    |
//| 473   | 1146 | R1 DATA |                                                                                                                                                    |
//| 473+E | 1146 | W0 DATA | @_SINT/CC/MAPR10NoCE1_ARA0 te=te:473 write(TCin1.9_V_5, C(TCin1.9_V_0)) @_SINT/CC/MAPR12NoCE1_ARB0 te=te:473 write(TCin1.9_V_5, C(TCin1.9_V_2))    |
//| 489   | 1146 | W1 DATA |                                                                                                                                                    |
//| 472   | 1147 | R0 DATA |                                                                                                                                                    |
//| 473   | 1147 | R1 DATA |                                                                                                                                                    |
//| 473+E | 1147 | W0 DATA | @_SINT/CC/MAPR10NoCE1_ARA0 te=te:473 write(TCin1.9_V_5, C(TCin1.9_V_0)) @_SINT/CC/MAPR12NoCE0_ARB0 te=te:473 write(TCin1.9_V_5, C(TCin1.9_V_2))    |
//| 490   | 1147 | W1 DATA |                                                                                                                                                    |
//| 472   | 1148 | R0 DATA |                                                                                                                                                    |
//| 473   | 1148 | R1 DATA |                                                                                                                                                    |
//| 473+E | 1148 | W0 DATA | @_SINT/CC/MAPR10NoCE1_ARA0 te=te:473 write(TCin1.9_V_5, C(TCin1.9_V_0)) TCi1._SPILL_256 te=te:473 scalarw(0)                                       |
//| 491   | 1148 | W1 DATA |                                                                                                                                                    |
//| 472   | 1149 | R0 DATA |                                                                                                                                                    |
//| 473   | 1149 | R1 DATA |                                                                                                                                                    |
//| 473+E | 1149 | W0 DATA | @_SINT/CC/MAPR10NoCE0_ARA0 te=te:473 write(TCin1.9_V_5, C(TCin1.9_V_0))  PLI:Eviction %u needed                                                    |
//| 492   | 1149 | W1 DATA |                                                                                                                                                    |
//| 472   | 1150 | R0 DATA |                                                                                                                                                    |
//| 473   | 1150 | R1 DATA |                                                                                                                                                    |
//| 473+E | 1150 | W0 DATA | @_SINT/CC/MAPR10NoCE0_ARA0 te=te:473 write(TCin1.9_V_5, C(TCin1.9_V_0)) @_SINT/CC/MAPR12NoCE3_ARB0 te=te:473 write(TCin1.9_V_5, C(TCin1.9_V_2))    |
//| 493   | 1150 | W1 DATA |                                                                                                                                                    |
//| 472   | 1151 | R0 DATA |                                                                                                                                                    |
//| 473   | 1151 | R1 DATA |                                                                                                                                                    |
//| 473+E | 1151 | W0 DATA | @_SINT/CC/MAPR10NoCE0_ARA0 te=te:473 write(TCin1.9_V_5, C(TCin1.9_V_0)) @_SINT/CC/MAPR12NoCE2_ARB0 te=te:473 write(TCin1.9_V_5, C(TCin1.9_V_2))    |
//| 494   | 1151 | W1 DATA |                                                                                                                                                    |
//| 472   | 1152 | R0 DATA |                                                                                                                                                    |
//| 473   | 1152 | R1 DATA |                                                                                                                                                    |
//| 473+E | 1152 | W0 DATA | @_SINT/CC/MAPR10NoCE0_ARA0 te=te:473 write(TCin1.9_V_5, C(TCin1.9_V_0)) @_SINT/CC/MAPR12NoCE1_ARB0 te=te:473 write(TCin1.9_V_5, C(TCin1.9_V_2))    |
//| 495   | 1152 | W1 DATA |                                                                                                                                                    |
//| 472   | 1153 | R0 DATA |                                                                                                                                                    |
//| 473   | 1153 | R1 DATA |                                                                                                                                                    |
//| 473+E | 1153 | W0 DATA | @_SINT/CC/MAPR10NoCE0_ARA0 te=te:473 write(TCin1.9_V_5, C(TCin1.9_V_0)) @_SINT/CC/MAPR12NoCE0_ARB0 te=te:473 write(TCin1.9_V_5, C(TCin1.9_V_2))    |
//| 496   | 1153 | W1 DATA |                                                                                                                                                    |
//| 472   | 1154 | R0 DATA |                                                                                                                                                    |
//| 473   | 1154 | R1 DATA |                                                                                                                                                    |
//| 473+E | 1154 | W0 DATA | @_SINT/CC/MAPR10NoCE0_ARA0 te=te:473 write(TCin1.9_V_5, C(TCin1.9_V_0)) TCi1._SPILL_256 te=te:473 scalarw(0)                                       |
//| 497   | 1154 | W1 DATA |                                                                                                                                                    |
//| 472   | 1155 | R0 DATA |                                                                                                                                                    |
//| 473   | 1155 | R1 DATA |                                                                                                                                                    |
//| 473+E | 1155 | W0 DATA | TCin1.9_V_1 te=te:473 scalarw(1+TCin1.9_V_1)  PLI:Eviction %u needed                                                                               |
//| 472   | 1156 | R0 DATA |                                                                                                                                                    |
//| 473   | 1156 | R1 DATA |                                                                                                                                                    |
//| 473+E | 1156 | W0 DATA | @_SINT/CC/MAPR12NoCE3_ARB0 te=te:473 write(TCin1.9_V_5, C(TCin1.9_V_2)) TCi1._SPILL_256 te=te:473 scalarw(0)                                       |
//| 498   | 1156 | W1 DATA |                                                                                                                                                    |
//| 472   | 1157 | R0 DATA |                                                                                                                                                    |
//| 473   | 1157 | R1 DATA |                                                                                                                                                    |
//| 473+E | 1157 | W0 DATA | @_SINT/CC/MAPR12NoCE2_ARB0 te=te:473 write(TCin1.9_V_5, C(TCin1.9_V_2)) TCi1._SPILL_256 te=te:473 scalarw(0)                                       |
//| 499   | 1157 | W1 DATA |                                                                                                                                                    |
//| 472   | 1158 | R0 DATA |                                                                                                                                                    |
//| 473   | 1158 | R1 DATA |                                                                                                                                                    |
//| 473+E | 1158 | W0 DATA | @_SINT/CC/MAPR12NoCE1_ARB0 te=te:473 write(TCin1.9_V_5, C(TCin1.9_V_2)) TCi1._SPILL_256 te=te:473 scalarw(0)                                       |
//| 500   | 1158 | W1 DATA |                                                                                                                                                    |
//| 472   | 1159 | R0 DATA |                                                                                                                                                    |
//| 473   | 1159 | R1 DATA |                                                                                                                                                    |
//| 473+E | 1159 | W0 DATA | @_SINT/CC/MAPR12NoCE0_ARB0 te=te:473 write(TCin1.9_V_5, C(TCin1.9_V_2)) TCi1._SPILL_256 te=te:473 scalarw(0)                                       |
//| 501   | 1159 | W1 DATA |                                                                                                                                                    |
//| 472   | 1160 | R0 DATA |                                                                                                                                                    |
//| 473   | 1160 | R1 DATA |                                                                                                                                                    |
//| 473+E | 1160 | W0 DATA | TTMT4Main_V_7 te=te:473 scalarw(S32'0I) TCi1._SPILL_256 te=te:473 scalarw(0)                                                                       |
//| 472   | 1161 | R0 DATA |                                                                                                                                                    |
//| 473   | 1161 | R1 DATA |                                                                                                                                                    |
//| 473+E | 1161 | W0 DATA | TCin1.9_V_4 te=te:473 scalarw(1+TCin1.9_V_4)                                                                                                       |
//*-------+------+---------+----------------------------------------------------------------------------------------------------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X95:"xpc10:95" 1162 :  major_start_pcl=502   edge_private_start/end=-1/-1 exec=502 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X95:"xpc10:95"
//res2: Thread=xpc10 state=X95:"xpc10:95"
//*-------+------+---------+----------------------------------------------*
//| pc    | eno  | Phaser  | Work                                         |
//*-------+------+---------+----------------------------------------------*
//| 502   | -    | R0 CTRL |                                              |
//| 502   | 1162 | R0 DATA |                                              |
//| 502+E | 1162 | W0 DATA | TCin1.9_V_1 te=te:502 scalarw(1+TCin1.9_V_1) |
//*-------+------+---------+----------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X96:"xpc10:96" 1189 :  major_start_pcl=503   edge_private_start/end=-1/-1 exec=503 (dend=0)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X96:"xpc10:96" 1188 :  major_start_pcl=503   edge_private_start/end=-1/-1 exec=503 (dend=0)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X96:"xpc10:96" 1187 :  major_start_pcl=503   edge_private_start/end=527/527 exec=503 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X96:"xpc10:96" 1186 :  major_start_pcl=503   edge_private_start/end=526/526 exec=503 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X96:"xpc10:96" 1185 :  major_start_pcl=503   edge_private_start/end=525/525 exec=503 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X96:"xpc10:96" 1184 :  major_start_pcl=503   edge_private_start/end=524/524 exec=503 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X96:"xpc10:96" 1183 :  major_start_pcl=503   edge_private_start/end=523/523 exec=503 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X96:"xpc10:96" 1182 :  major_start_pcl=503   edge_private_start/end=522/522 exec=503 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X96:"xpc10:96" 1181 :  major_start_pcl=503   edge_private_start/end=521/521 exec=503 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X96:"xpc10:96" 1180 :  major_start_pcl=503   edge_private_start/end=520/520 exec=503 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X96:"xpc10:96" 1179 :  major_start_pcl=503   edge_private_start/end=519/519 exec=503 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X96:"xpc10:96" 1178 :  major_start_pcl=503   edge_private_start/end=518/518 exec=503 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X96:"xpc10:96" 1177 :  major_start_pcl=503   edge_private_start/end=517/517 exec=503 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X96:"xpc10:96" 1176 :  major_start_pcl=503   edge_private_start/end=516/516 exec=503 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X96:"xpc10:96" 1175 :  major_start_pcl=503   edge_private_start/end=515/515 exec=503 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X96:"xpc10:96" 1174 :  major_start_pcl=503   edge_private_start/end=514/514 exec=503 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X96:"xpc10:96" 1173 :  major_start_pcl=503   edge_private_start/end=513/513 exec=503 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X96:"xpc10:96" 1172 :  major_start_pcl=503   edge_private_start/end=512/512 exec=503 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X96:"xpc10:96" 1171 :  major_start_pcl=503   edge_private_start/end=511/511 exec=503 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X96:"xpc10:96" 1170 :  major_start_pcl=503   edge_private_start/end=510/510 exec=503 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X96:"xpc10:96" 1169 :  major_start_pcl=503   edge_private_start/end=509/509 exec=503 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X96:"xpc10:96" 1168 :  major_start_pcl=503   edge_private_start/end=508/508 exec=503 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X96:"xpc10:96" 1167 :  major_start_pcl=503   edge_private_start/end=507/507 exec=503 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X96:"xpc10:96" 1166 :  major_start_pcl=503   edge_private_start/end=506/506 exec=503 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X96:"xpc10:96" 1165 :  major_start_pcl=503   edge_private_start/end=505/505 exec=503 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X96:"xpc10:96" 1164 :  major_start_pcl=503   edge_private_start/end=504/504 exec=503 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X96:"xpc10:96" 1163 :  major_start_pcl=503   edge_private_start/end=-1/-1 exec=503 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X96:"xpc10:96"
//res2: Thread=xpc10 state=X96:"xpc10:96"
//*-------+------+---------+-------------------------------------------------------------------------------------------------------------------------------------------------*
//| pc    | eno  | Phaser  | Work                                                                                                                                            |
//*-------+------+---------+-------------------------------------------------------------------------------------------------------------------------------------------------*
//| 503   | -    | R0 CTRL |                                                                                                                                                 |
//| 503   | 1163 | R0 DATA |                                                                                                                                                 |
//| 503+E | 1163 | W0 DATA | TCin1.9_V_1 te=te:503 scalarw(1+TCin1.9_V_1) @_SINT/CC/SCALbx24_stats_insert_probes te=te:503 scalarw(E13)  PLI:Eviction %u needed              |
//| 503   | 1164 | R0 DATA |                                                                                                                                                 |
//| 503+E | 1164 | W0 DATA | @_SINT/CC/MAPR10NoCE3_ARA0 te=te:503 write(TCin1.9_V_5, C(TCin1.9_V_0)) @_SINT/CC/MAPR12NoCE3_ARB0 te=te:503 write(TCin1.9_V_5, C(TCin1.9_V_2)) |
//| 504   | 1164 | W1 DATA |                                                                                                                                                 |
//| 503   | 1165 | R0 DATA |                                                                                                                                                 |
//| 503+E | 1165 | W0 DATA | @_SINT/CC/MAPR10NoCE3_ARA0 te=te:503 write(TCin1.9_V_5, C(TCin1.9_V_0)) @_SINT/CC/MAPR12NoCE2_ARB0 te=te:503 write(TCin1.9_V_5, C(TCin1.9_V_2)) |
//| 505   | 1165 | W1 DATA |                                                                                                                                                 |
//| 503   | 1166 | R0 DATA |                                                                                                                                                 |
//| 503+E | 1166 | W0 DATA | @_SINT/CC/MAPR10NoCE3_ARA0 te=te:503 write(TCin1.9_V_5, C(TCin1.9_V_0)) @_SINT/CC/MAPR12NoCE1_ARB0 te=te:503 write(TCin1.9_V_5, C(TCin1.9_V_2)) |
//| 506   | 1166 | W1 DATA |                                                                                                                                                 |
//| 503   | 1167 | R0 DATA |                                                                                                                                                 |
//| 503+E | 1167 | W0 DATA | @_SINT/CC/MAPR10NoCE3_ARA0 te=te:503 write(TCin1.9_V_5, C(TCin1.9_V_0)) @_SINT/CC/MAPR12NoCE0_ARB0 te=te:503 write(TCin1.9_V_5, C(TCin1.9_V_2)) |
//| 507   | 1167 | W1 DATA |                                                                                                                                                 |
//| 503   | 1168 | R0 DATA |                                                                                                                                                 |
//| 503+E | 1168 | W0 DATA | @_SINT/CC/MAPR10NoCE3_ARA0 te=te:503 write(TCin1.9_V_5, C(TCin1.9_V_0)) TCi1._SPILL_256 te=te:503 scalarw(0)                                    |
//| 508   | 1168 | W1 DATA |                                                                                                                                                 |
//| 503   | 1169 | R0 DATA |                                                                                                                                                 |
//| 503+E | 1169 | W0 DATA | @_SINT/CC/MAPR10NoCE2_ARA0 te=te:503 write(TCin1.9_V_5, C(TCin1.9_V_0)) @_SINT/CC/MAPR12NoCE3_ARB0 te=te:503 write(TCin1.9_V_5, C(TCin1.9_V_2)) |
//| 509   | 1169 | W1 DATA |                                                                                                                                                 |
//| 503   | 1170 | R0 DATA |                                                                                                                                                 |
//| 503+E | 1170 | W0 DATA | @_SINT/CC/MAPR10NoCE2_ARA0 te=te:503 write(TCin1.9_V_5, C(TCin1.9_V_0)) @_SINT/CC/MAPR12NoCE2_ARB0 te=te:503 write(TCin1.9_V_5, C(TCin1.9_V_2)) |
//| 510   | 1170 | W1 DATA |                                                                                                                                                 |
//| 503   | 1171 | R0 DATA |                                                                                                                                                 |
//| 503+E | 1171 | W0 DATA | @_SINT/CC/MAPR10NoCE2_ARA0 te=te:503 write(TCin1.9_V_5, C(TCin1.9_V_0)) @_SINT/CC/MAPR12NoCE1_ARB0 te=te:503 write(TCin1.9_V_5, C(TCin1.9_V_2)) |
//| 511   | 1171 | W1 DATA |                                                                                                                                                 |
//| 503   | 1172 | R0 DATA |                                                                                                                                                 |
//| 503+E | 1172 | W0 DATA | @_SINT/CC/MAPR10NoCE2_ARA0 te=te:503 write(TCin1.9_V_5, C(TCin1.9_V_0)) @_SINT/CC/MAPR12NoCE0_ARB0 te=te:503 write(TCin1.9_V_5, C(TCin1.9_V_2)) |
//| 512   | 1172 | W1 DATA |                                                                                                                                                 |
//| 503   | 1173 | R0 DATA |                                                                                                                                                 |
//| 503+E | 1173 | W0 DATA | @_SINT/CC/MAPR10NoCE2_ARA0 te=te:503 write(TCin1.9_V_5, C(TCin1.9_V_0)) TCi1._SPILL_256 te=te:503 scalarw(0)                                    |
//| 513   | 1173 | W1 DATA |                                                                                                                                                 |
//| 503   | 1174 | R0 DATA |                                                                                                                                                 |
//| 503+E | 1174 | W0 DATA | @_SINT/CC/MAPR10NoCE1_ARA0 te=te:503 write(TCin1.9_V_5, C(TCin1.9_V_0)) @_SINT/CC/MAPR12NoCE3_ARB0 te=te:503 write(TCin1.9_V_5, C(TCin1.9_V_2)) |
//| 514   | 1174 | W1 DATA |                                                                                                                                                 |
//| 503   | 1175 | R0 DATA |                                                                                                                                                 |
//| 503+E | 1175 | W0 DATA | @_SINT/CC/MAPR10NoCE1_ARA0 te=te:503 write(TCin1.9_V_5, C(TCin1.9_V_0)) @_SINT/CC/MAPR12NoCE2_ARB0 te=te:503 write(TCin1.9_V_5, C(TCin1.9_V_2)) |
//| 515   | 1175 | W1 DATA |                                                                                                                                                 |
//| 503   | 1176 | R0 DATA |                                                                                                                                                 |
//| 503+E | 1176 | W0 DATA | @_SINT/CC/MAPR10NoCE1_ARA0 te=te:503 write(TCin1.9_V_5, C(TCin1.9_V_0)) @_SINT/CC/MAPR12NoCE1_ARB0 te=te:503 write(TCin1.9_V_5, C(TCin1.9_V_2)) |
//| 516   | 1176 | W1 DATA |                                                                                                                                                 |
//| 503   | 1177 | R0 DATA |                                                                                                                                                 |
//| 503+E | 1177 | W0 DATA | @_SINT/CC/MAPR10NoCE1_ARA0 te=te:503 write(TCin1.9_V_5, C(TCin1.9_V_0)) @_SINT/CC/MAPR12NoCE0_ARB0 te=te:503 write(TCin1.9_V_5, C(TCin1.9_V_2)) |
//| 517   | 1177 | W1 DATA |                                                                                                                                                 |
//| 503   | 1178 | R0 DATA |                                                                                                                                                 |
//| 503+E | 1178 | W0 DATA | @_SINT/CC/MAPR10NoCE1_ARA0 te=te:503 write(TCin1.9_V_5, C(TCin1.9_V_0)) TCi1._SPILL_256 te=te:503 scalarw(0)                                    |
//| 518   | 1178 | W1 DATA |                                                                                                                                                 |
//| 503   | 1179 | R0 DATA |                                                                                                                                                 |
//| 503+E | 1179 | W0 DATA | @_SINT/CC/MAPR10NoCE0_ARA0 te=te:503 write(TCin1.9_V_5, C(TCin1.9_V_0)) @_SINT/CC/MAPR12NoCE3_ARB0 te=te:503 write(TCin1.9_V_5, C(TCin1.9_V_2)) |
//| 519   | 1179 | W1 DATA |                                                                                                                                                 |
//| 503   | 1180 | R0 DATA |                                                                                                                                                 |
//| 503+E | 1180 | W0 DATA | @_SINT/CC/MAPR10NoCE0_ARA0 te=te:503 write(TCin1.9_V_5, C(TCin1.9_V_0)) @_SINT/CC/MAPR12NoCE2_ARB0 te=te:503 write(TCin1.9_V_5, C(TCin1.9_V_2)) |
//| 520   | 1180 | W1 DATA |                                                                                                                                                 |
//| 503   | 1181 | R0 DATA |                                                                                                                                                 |
//| 503+E | 1181 | W0 DATA | @_SINT/CC/MAPR10NoCE0_ARA0 te=te:503 write(TCin1.9_V_5, C(TCin1.9_V_0)) @_SINT/CC/MAPR12NoCE1_ARB0 te=te:503 write(TCin1.9_V_5, C(TCin1.9_V_2)) |
//| 521   | 1181 | W1 DATA |                                                                                                                                                 |
//| 503   | 1182 | R0 DATA |                                                                                                                                                 |
//| 503+E | 1182 | W0 DATA | @_SINT/CC/MAPR10NoCE0_ARA0 te=te:503 write(TCin1.9_V_5, C(TCin1.9_V_0)) @_SINT/CC/MAPR12NoCE0_ARB0 te=te:503 write(TCin1.9_V_5, C(TCin1.9_V_2)) |
//| 522   | 1182 | W1 DATA |                                                                                                                                                 |
//| 503   | 1183 | R0 DATA |                                                                                                                                                 |
//| 503+E | 1183 | W0 DATA | @_SINT/CC/MAPR10NoCE0_ARA0 te=te:503 write(TCin1.9_V_5, C(TCin1.9_V_0)) TCi1._SPILL_256 te=te:503 scalarw(0)                                    |
//| 523   | 1183 | W1 DATA |                                                                                                                                                 |
//| 503   | 1184 | R0 DATA |                                                                                                                                                 |
//| 503+E | 1184 | W0 DATA | @_SINT/CC/MAPR12NoCE3_ARB0 te=te:503 write(TCin1.9_V_5, C(TCin1.9_V_2)) TCi1._SPILL_256 te=te:503 scalarw(0)                                    |
//| 524   | 1184 | W1 DATA |                                                                                                                                                 |
//| 503   | 1185 | R0 DATA |                                                                                                                                                 |
//| 503+E | 1185 | W0 DATA | @_SINT/CC/MAPR12NoCE2_ARB0 te=te:503 write(TCin1.9_V_5, C(TCin1.9_V_2)) TCi1._SPILL_256 te=te:503 scalarw(0)                                    |
//| 525   | 1185 | W1 DATA |                                                                                                                                                 |
//| 503   | 1186 | R0 DATA |                                                                                                                                                 |
//| 503+E | 1186 | W0 DATA | @_SINT/CC/MAPR12NoCE1_ARB0 te=te:503 write(TCin1.9_V_5, C(TCin1.9_V_2)) TCi1._SPILL_256 te=te:503 scalarw(0)                                    |
//| 526   | 1186 | W1 DATA |                                                                                                                                                 |
//| 503   | 1187 | R0 DATA |                                                                                                                                                 |
//| 503+E | 1187 | W0 DATA | @_SINT/CC/MAPR12NoCE0_ARB0 te=te:503 write(TCin1.9_V_5, C(TCin1.9_V_2)) TCi1._SPILL_256 te=te:503 scalarw(0)                                    |
//| 527   | 1187 | W1 DATA |                                                                                                                                                 |
//| 503   | 1188 | R0 DATA |                                                                                                                                                 |
//| 503+E | 1188 | W0 DATA | TTMT4Main_V_7 te=te:503 scalarw(S32'0I) TCi1._SPILL_256 te=te:503 scalarw(0)                                                                    |
//| 503   | 1189 | R0 DATA |                                                                                                                                                 |
//| 503+E | 1189 | W0 DATA | TCin1.9_V_1 te=te:503 scalarw(1+TCin1.9_V_1) @_SINT/CC/SCALbx24_stats_insert_probes te=te:503 scalarw(E13)  PLI:Eviction %u needed              |
//*-------+------+---------+-------------------------------------------------------------------------------------------------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X97:"xpc10:97" 1193 :  major_start_pcl=528   edge_private_start/end=-1/-1 exec=528 (dend=0)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X97:"xpc10:97" 1192 :  major_start_pcl=528   edge_private_start/end=531/531 exec=528 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X97:"xpc10:97" 1191 :  major_start_pcl=528   edge_private_start/end=530/530 exec=528 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X97:"xpc10:97" 1190 :  major_start_pcl=528   edge_private_start/end=529/529 exec=528 (dend=1)
//Simple greedy schedule for res2: Thread=xpc10 state=X97:"xpc10:97"
//res2: Thread=xpc10 state=X97:"xpc10:97"
//*-------+------+---------+------------------------------------------------------------------------------------------------------------*
//| pc    | eno  | Phaser  | Work                                                                                                       |
//*-------+------+---------+------------------------------------------------------------------------------------------------------------*
//| 528   | -    | R0 CTRL |                                                                                                            |
//| 528   | 1190 | R0 DATA |                                                                                                            |
//| 528+E | 1190 | W0 DATA | TCCl0.12_V_1 te=te:528 scalarw(1+TCCl0.12_V_1) @_SINT/CC/MAPR10NoCE2_ARA0 te=te:528 write(TCCl0.12_V_0, 0) |
//| 529   | 1190 | W1 DATA |                                                                                                            |
//| 528   | 1191 | R0 DATA |                                                                                                            |
//| 528+E | 1191 | W0 DATA | TCCl0.12_V_1 te=te:528 scalarw(1+TCCl0.12_V_1) @_SINT/CC/MAPR10NoCE1_ARA0 te=te:528 write(TCCl0.12_V_0, 0) |
//| 530   | 1191 | W1 DATA |                                                                                                            |
//| 528   | 1192 | R0 DATA |                                                                                                            |
//| 528+E | 1192 | W0 DATA | TCCl0.12_V_1 te=te:528 scalarw(1+TCCl0.12_V_1) @_SINT/CC/MAPR10NoCE0_ARA0 te=te:528 write(TCCl0.12_V_0, 0) |
//| 531   | 1192 | W1 DATA |                                                                                                            |
//| 528   | 1193 | R0 DATA |                                                                                                            |
//| 528+E | 1193 | W0 DATA | TCCl0.12_V_1 te=te:528 scalarw(1+TCCl0.12_V_1)                                                             |
//*-------+------+---------+------------------------------------------------------------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X98:"xpc10:98" 1195 :  major_start_pcl=532   edge_private_start/end=-1/-1 exec=532 (dend=0)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X98:"xpc10:98" 1194 :  major_start_pcl=532   edge_private_start/end=533/533 exec=532 (dend=1)
//Simple greedy schedule for res2: Thread=xpc10 state=X98:"xpc10:98"
//res2: Thread=xpc10 state=X98:"xpc10:98"
//*-------+------+---------+--------------------------------------------------------------------------------------------------------------------------------*
//| pc    | eno  | Phaser  | Work                                                                                                                           |
//*-------+------+---------+--------------------------------------------------------------------------------------------------------------------------------*
//| 532   | -    | R0 CTRL |                                                                                                                                |
//| 532   | 1194 | R0 DATA |                                                                                                                                |
//| 532+E | 1194 | W0 DATA | TCCl0.12_V_1 te=te:532 scalarw(1+TCCl0.12_V_1) @_SINT/CC/MAPR10NoCE3_ARA0 te=te:532 write(TCCl0.12_V_0, 0) @_SINT/CC/MAPR10No\ |
//|       |      |         | CE2_ARA0 te=te:532 write(TCCl0.12_V_0, 0) @_SINT/CC/MAPR10NoCE1_ARA0 te=te:532 write(TCCl0.12_V_0, 0) @_SINT/CC/MAPR10NoCE0_A\ |
//|       |      |         | RA0 te=te:532 write(TCCl0.12_V_0, 0)                                                                                           |
//| 533   | 1194 | W1 DATA |                                                                                                                                |
//| 532   | 1195 | R0 DATA |                                                                                                                                |
//| 532+E | 1195 | W0 DATA | TCCl0.12_V_0 te=te:532 scalarw(1+TCCl0.12_V_0)                                                                                 |
//*-------+------+---------+--------------------------------------------------------------------------------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X99:"xpc10:99" 1198 :  major_start_pcl=534   edge_private_start/end=-1/-1 exec=534 (dend=0)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X99:"xpc10:99" 1197 :  major_start_pcl=534   edge_private_start/end=536/536 exec=534 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X99:"xpc10:99" 1196 :  major_start_pcl=534   edge_private_start/end=535/535 exec=534 (dend=1)
//Simple greedy schedule for res2: Thread=xpc10 state=X99:"xpc10:99"
//res2: Thread=xpc10 state=X99:"xpc10:99"
//*-------+------+---------+------------------------------------------------------------------------------------------------------------*
//| pc    | eno  | Phaser  | Work                                                                                                       |
//*-------+------+---------+------------------------------------------------------------------------------------------------------------*
//| 534   | -    | R0 CTRL |                                                                                                            |
//| 534   | 1196 | R0 DATA |                                                                                                            |
//| 534+E | 1196 | W0 DATA | TCCl0.12_V_1 te=te:534 scalarw(1+TCCl0.12_V_1) @_SINT/CC/MAPR10NoCE1_ARA0 te=te:534 write(TCCl0.12_V_0, 0) |
//| 535   | 1196 | W1 DATA |                                                                                                            |
//| 534   | 1197 | R0 DATA |                                                                                                            |
//| 534+E | 1197 | W0 DATA | TCCl0.12_V_1 te=te:534 scalarw(1+TCCl0.12_V_1) @_SINT/CC/MAPR10NoCE0_ARA0 te=te:534 write(TCCl0.12_V_0, 0) |
//| 536   | 1197 | W1 DATA |                                                                                                            |
//| 534   | 1198 | R0 DATA |                                                                                                            |
//| 534+E | 1198 | W0 DATA | TCCl0.12_V_1 te=te:534 scalarw(1+TCCl0.12_V_1)                                                             |
//*-------+------+---------+------------------------------------------------------------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X100:"xpc10:100" 1200 :  major_start_pcl=537   edge_private_start/end=-1/-1 exec=537 (dend=0)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X100:"xpc10:100" 1199 :  major_start_pcl=537   edge_private_start/end=538/538 exec=537 (dend=1)
//Simple greedy schedule for res2: Thread=xpc10 state=X100:"xpc10:100"
//res2: Thread=xpc10 state=X100:"xpc10:100"
//*-------+------+---------+------------------------------------------------------------------------------------------------------------*
//| pc    | eno  | Phaser  | Work                                                                                                       |
//*-------+------+---------+------------------------------------------------------------------------------------------------------------*
//| 537   | -    | R0 CTRL |                                                                                                            |
//| 537   | 1199 | R0 DATA |                                                                                                            |
//| 537+E | 1199 | W0 DATA | TCCl0.12_V_1 te=te:537 scalarw(1+TCCl0.12_V_1) @_SINT/CC/MAPR10NoCE0_ARA0 te=te:537 write(TCCl0.12_V_0, 0) |
//| 538   | 1199 | W1 DATA |                                                                                                            |
//| 537   | 1200 | R0 DATA |                                                                                                            |
//| 537+E | 1200 | W0 DATA | TCCl0.12_V_1 te=te:537 scalarw(1+TCCl0.12_V_1)                                                             |
//*-------+------+---------+------------------------------------------------------------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X101:"xpc10:101" 1201 :  major_start_pcl=539   edge_private_start/end=-1/-1 exec=539 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X101:"xpc10:101"
//res2: Thread=xpc10 state=X101:"xpc10:101"
//*-------+------+---------+------------------------------------------------*
//| pc    | eno  | Phaser  | Work                                           |
//*-------+------+---------+------------------------------------------------*
//| 539   | -    | R0 CTRL |                                                |
//| 539   | 1201 | R0 DATA |                                                |
//| 539+E | 1201 | W0 DATA | TCCl0.12_V_1 te=te:539 scalarw(1+TCCl0.12_V_1) |
//*-------+------+---------+------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X102:"xpc10:102" 1205 :  major_start_pcl=540   edge_private_start/end=-1/-1 exec=540 (dend=0)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X102:"xpc10:102" 1204 :  major_start_pcl=540   edge_private_start/end=543/543 exec=540 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X102:"xpc10:102" 1203 :  major_start_pcl=540   edge_private_start/end=542/542 exec=540 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X102:"xpc10:102" 1202 :  major_start_pcl=540   edge_private_start/end=541/541 exec=540 (dend=1)
//Simple greedy schedule for res2: Thread=xpc10 state=X102:"xpc10:102"
//res2: Thread=xpc10 state=X102:"xpc10:102"
//*-------+------+---------+------------------------------------------------------------------------------------*
//| pc    | eno  | Phaser  | Work                                                                               |
//*-------+------+---------+------------------------------------------------------------------------------------*
//| 540   | -    | R0 CTRL |                                                                                    |
//| 540   | 1202 | R0 DATA |                                                                                    |
//| 540+E | 1202 | W0 DATA | TCCl0.12_V_1 te=te:540 scalarw(4) @_SINT/CC/MAPR10NoCE2_ARA0 te=te:540 write(0, 0) |
//| 541   | 1202 | W1 DATA |                                                                                    |
//| 540   | 1203 | R0 DATA |                                                                                    |
//| 540+E | 1203 | W0 DATA | TCCl0.12_V_1 te=te:540 scalarw(4) @_SINT/CC/MAPR10NoCE1_ARA0 te=te:540 write(0, 0) |
//| 542   | 1203 | W1 DATA |                                                                                    |
//| 540   | 1204 | R0 DATA |                                                                                    |
//| 540+E | 1204 | W0 DATA | TCCl0.12_V_1 te=te:540 scalarw(4) @_SINT/CC/MAPR10NoCE0_ARA0 te=te:540 write(0, 0) |
//| 543   | 1204 | W1 DATA |                                                                                    |
//| 540   | 1205 | R0 DATA |                                                                                    |
//| 540+E | 1205 | W0 DATA | TCCl0.12_V_1 te=te:540 scalarw(4) TCCl0.12_V_0 te=te:540 scalarw(1+TCCl0.12_V_0)   |
//*-------+------+---------+------------------------------------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X103:"xpc10:103" 1208 :  major_start_pcl=544   edge_private_start/end=-1/-1 exec=544 (dend=0)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X103:"xpc10:103" 1207 :  major_start_pcl=544   edge_private_start/end=546/546 exec=544 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X103:"xpc10:103" 1206 :  major_start_pcl=544   edge_private_start/end=545/545 exec=544 (dend=1)
//Simple greedy schedule for res2: Thread=xpc10 state=X103:"xpc10:103"
//res2: Thread=xpc10 state=X103:"xpc10:103"
//*-------+------+---------+------------------------------------------------------------------------------------*
//| pc    | eno  | Phaser  | Work                                                                               |
//*-------+------+---------+------------------------------------------------------------------------------------*
//| 544   | -    | R0 CTRL |                                                                                    |
//| 544   | 1206 | R0 DATA |                                                                                    |
//| 544+E | 1206 | W0 DATA | TCCl0.12_V_1 te=te:544 scalarw(4) @_SINT/CC/MAPR10NoCE1_ARA0 te=te:544 write(0, 0) |
//| 545   | 1206 | W1 DATA |                                                                                    |
//| 544   | 1207 | R0 DATA |                                                                                    |
//| 544+E | 1207 | W0 DATA | TCCl0.12_V_1 te=te:544 scalarw(4) @_SINT/CC/MAPR10NoCE0_ARA0 te=te:544 write(0, 0) |
//| 546   | 1207 | W1 DATA |                                                                                    |
//| 544   | 1208 | R0 DATA |                                                                                    |
//| 544+E | 1208 | W0 DATA | TCCl0.12_V_1 te=te:544 scalarw(4) TCCl0.12_V_0 te=te:544 scalarw(1+TCCl0.12_V_0)   |
//*-------+------+---------+------------------------------------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X104:"xpc10:104" 1210 :  major_start_pcl=547   edge_private_start/end=-1/-1 exec=547 (dend=0)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X104:"xpc10:104" 1209 :  major_start_pcl=547   edge_private_start/end=548/548 exec=547 (dend=1)
//Simple greedy schedule for res2: Thread=xpc10 state=X104:"xpc10:104"
//res2: Thread=xpc10 state=X104:"xpc10:104"
//*-------+------+---------+------------------------------------------------------------------------------------*
//| pc    | eno  | Phaser  | Work                                                                               |
//*-------+------+---------+------------------------------------------------------------------------------------*
//| 547   | -    | R0 CTRL |                                                                                    |
//| 547   | 1209 | R0 DATA |                                                                                    |
//| 547+E | 1209 | W0 DATA | TCCl0.12_V_1 te=te:547 scalarw(4) @_SINT/CC/MAPR10NoCE0_ARA0 te=te:547 write(0, 0) |
//| 548   | 1209 | W1 DATA |                                                                                    |
//| 547   | 1210 | R0 DATA |                                                                                    |
//| 547+E | 1210 | W0 DATA | TCCl0.12_V_1 te=te:547 scalarw(4) TCCl0.12_V_0 te=te:547 scalarw(1+TCCl0.12_V_0)   |
//*-------+------+---------+------------------------------------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X105:"xpc10:105" 1211 :  major_start_pcl=549   edge_private_start/end=-1/-1 exec=549 (dend=0)
//Simple greedy schedule for res2: Thread=xpc10 state=X105:"xpc10:105"
//res2: Thread=xpc10 state=X105:"xpc10:105"
//*-------+------+---------+----------------------------------------------------------------------------------*
//| pc    | eno  | Phaser  | Work                                                                             |
//*-------+------+---------+----------------------------------------------------------------------------------*
//| 549   | -    | R0 CTRL |                                                                                  |
//| 549   | 1211 | R0 DATA |                                                                                  |
//| 549+E | 1211 | W0 DATA | TCCl0.12_V_1 te=te:549 scalarw(4) TCCl0.12_V_0 te=te:549 scalarw(1+TCCl0.12_V_0) |
//*-------+------+---------+----------------------------------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X106:"xpc10:106" 1219 :  major_start_pcl=550   edge_private_start/end=-1/-1 exec=550 (dend=0)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X106:"xpc10:106" 1218 :  major_start_pcl=550   edge_private_start/end=557/557 exec=550 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X106:"xpc10:106" 1217 :  major_start_pcl=550   edge_private_start/end=556/556 exec=550 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X106:"xpc10:106" 1216 :  major_start_pcl=550   edge_private_start/end=555/555 exec=550 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X106:"xpc10:106" 1215 :  major_start_pcl=550   edge_private_start/end=554/554 exec=550 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X106:"xpc10:106" 1214 :  major_start_pcl=550   edge_private_start/end=553/553 exec=550 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X106:"xpc10:106" 1213 :  major_start_pcl=550   edge_private_start/end=552/552 exec=550 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X106:"xpc10:106" 1212 :  major_start_pcl=550   edge_private_start/end=551/551 exec=550 (dend=1)
//Simple greedy schedule for res2: Thread=xpc10 state=X106:"xpc10:106"
//res2: Thread=xpc10 state=X106:"xpc10:106"
//*-------+------+---------+------------------------------------------------------------------------------------*
//| pc    | eno  | Phaser  | Work                                                                               |
//*-------+------+---------+------------------------------------------------------------------------------------*
//| 550   | -    | R0 CTRL |                                                                                    |
//| 550   | 1212 | R0 DATA |                                                                                    |
//| 550+E | 1212 | W0 DATA | TCCl0.12_V_1 te=te:550 scalarw(3) @_SINT/CC/MAPR10NoCE2_ARA0 te=te:550 write(0, 0) |
//| 551   | 1212 | W1 DATA |                                                                                    |
//| 550   | 1213 | R0 DATA |                                                                                    |
//| 550+E | 1213 | W0 DATA | TCCl0.12_V_1 te=te:550 scalarw(3) @_SINT/CC/MAPR10NoCE1_ARA0 te=te:550 write(0, 0) |
//| 552   | 1213 | W1 DATA |                                                                                    |
//| 550   | 1214 | R0 DATA |                                                                                    |
//| 550+E | 1214 | W0 DATA | TCCl0.12_V_1 te=te:550 scalarw(3) @_SINT/CC/MAPR10NoCE0_ARA0 te=te:550 write(0, 0) |
//| 553   | 1214 | W1 DATA |                                                                                    |
//| 550   | 1215 | R0 DATA |                                                                                    |
//| 550+E | 1215 | W0 DATA | TCCl0.12_V_1 te=te:550 scalarw(3) @_SINT/CC/MAPR10NoCE3_ARA0 te=te:550 write(0, 0) |
//| 554   | 1215 | W1 DATA |                                                                                    |
//| 550   | 1216 | R0 DATA |                                                                                    |
//| 550+E | 1216 | W0 DATA | TCCl0.12_V_1 te=te:550 scalarw(3) @_SINT/CC/MAPR10NoCE2_ARA0 te=te:550 write(0, 0) |
//| 555   | 1216 | W1 DATA |                                                                                    |
//| 550   | 1217 | R0 DATA |                                                                                    |
//| 550+E | 1217 | W0 DATA | TCCl0.12_V_1 te=te:550 scalarw(3) @_SINT/CC/MAPR10NoCE1_ARA0 te=te:550 write(0, 0) |
//| 556   | 1217 | W1 DATA |                                                                                    |
//| 550   | 1218 | R0 DATA |                                                                                    |
//| 550+E | 1218 | W0 DATA | TCCl0.12_V_1 te=te:550 scalarw(3) @_SINT/CC/MAPR10NoCE0_ARA0 te=te:550 write(0, 0) |
//| 557   | 1218 | W1 DATA |                                                                                    |
//| 550   | 1219 | R0 DATA |                                                                                    |
//| 550+E | 1219 | W0 DATA | TCCl0.12_V_1 te=te:550 scalarw(4) TCCl0.12_V_0 te=te:550 scalarw(1+TCCl0.12_V_0)   |
//*-------+------+---------+------------------------------------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X107:"xpc10:107" 1226 :  major_start_pcl=558   edge_private_start/end=-1/-1 exec=558 (dend=0)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X107:"xpc10:107" 1225 :  major_start_pcl=558   edge_private_start/end=564/564 exec=558 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X107:"xpc10:107" 1224 :  major_start_pcl=558   edge_private_start/end=563/563 exec=558 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X107:"xpc10:107" 1223 :  major_start_pcl=558   edge_private_start/end=562/562 exec=558 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X107:"xpc10:107" 1222 :  major_start_pcl=558   edge_private_start/end=561/561 exec=558 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X107:"xpc10:107" 1221 :  major_start_pcl=558   edge_private_start/end=560/560 exec=558 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X107:"xpc10:107" 1220 :  major_start_pcl=558   edge_private_start/end=559/559 exec=558 (dend=1)
//Simple greedy schedule for res2: Thread=xpc10 state=X107:"xpc10:107"
//res2: Thread=xpc10 state=X107:"xpc10:107"
//*-------+------+---------+------------------------------------------------------------------------------------*
//| pc    | eno  | Phaser  | Work                                                                               |
//*-------+------+---------+------------------------------------------------------------------------------------*
//| 558   | -    | R0 CTRL |                                                                                    |
//| 558   | 1220 | R0 DATA |                                                                                    |
//| 558+E | 1220 | W0 DATA | TCCl0.12_V_1 te=te:558 scalarw(3) @_SINT/CC/MAPR10NoCE1_ARA0 te=te:558 write(0, 0) |
//| 559   | 1220 | W1 DATA |                                                                                    |
//| 558   | 1221 | R0 DATA |                                                                                    |
//| 558+E | 1221 | W0 DATA | TCCl0.12_V_1 te=te:558 scalarw(3) @_SINT/CC/MAPR10NoCE0_ARA0 te=te:558 write(0, 0) |
//| 560   | 1221 | W1 DATA |                                                                                    |
//| 558   | 1222 | R0 DATA |                                                                                    |
//| 558+E | 1222 | W0 DATA | TCCl0.12_V_1 te=te:558 scalarw(3) @_SINT/CC/MAPR10NoCE3_ARA0 te=te:558 write(0, 0) |
//| 561   | 1222 | W1 DATA |                                                                                    |
//| 558   | 1223 | R0 DATA |                                                                                    |
//| 558+E | 1223 | W0 DATA | TCCl0.12_V_1 te=te:558 scalarw(3) @_SINT/CC/MAPR10NoCE2_ARA0 te=te:558 write(0, 0) |
//| 562   | 1223 | W1 DATA |                                                                                    |
//| 558   | 1224 | R0 DATA |                                                                                    |
//| 558+E | 1224 | W0 DATA | TCCl0.12_V_1 te=te:558 scalarw(3) @_SINT/CC/MAPR10NoCE1_ARA0 te=te:558 write(0, 0) |
//| 563   | 1224 | W1 DATA |                                                                                    |
//| 558   | 1225 | R0 DATA |                                                                                    |
//| 558+E | 1225 | W0 DATA | TCCl0.12_V_1 te=te:558 scalarw(3) @_SINT/CC/MAPR10NoCE0_ARA0 te=te:558 write(0, 0) |
//| 564   | 1225 | W1 DATA |                                                                                    |
//| 558   | 1226 | R0 DATA |                                                                                    |
//| 558+E | 1226 | W0 DATA | TCCl0.12_V_1 te=te:558 scalarw(4) TCCl0.12_V_0 te=te:558 scalarw(1+TCCl0.12_V_0)   |
//*-------+------+---------+------------------------------------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X108:"xpc10:108" 1232 :  major_start_pcl=565   edge_private_start/end=-1/-1 exec=565 (dend=0)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X108:"xpc10:108" 1231 :  major_start_pcl=565   edge_private_start/end=570/570 exec=565 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X108:"xpc10:108" 1230 :  major_start_pcl=565   edge_private_start/end=569/569 exec=565 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X108:"xpc10:108" 1229 :  major_start_pcl=565   edge_private_start/end=568/568 exec=565 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X108:"xpc10:108" 1228 :  major_start_pcl=565   edge_private_start/end=567/567 exec=565 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X108:"xpc10:108" 1227 :  major_start_pcl=565   edge_private_start/end=566/566 exec=565 (dend=1)
//Simple greedy schedule for res2: Thread=xpc10 state=X108:"xpc10:108"
//res2: Thread=xpc10 state=X108:"xpc10:108"
//*-------+------+---------+------------------------------------------------------------------------------------*
//| pc    | eno  | Phaser  | Work                                                                               |
//*-------+------+---------+------------------------------------------------------------------------------------*
//| 565   | -    | R0 CTRL |                                                                                    |
//| 565   | 1227 | R0 DATA |                                                                                    |
//| 565+E | 1227 | W0 DATA | TCCl0.12_V_1 te=te:565 scalarw(3) @_SINT/CC/MAPR10NoCE0_ARA0 te=te:565 write(0, 0) |
//| 566   | 1227 | W1 DATA |                                                                                    |
//| 565   | 1228 | R0 DATA |                                                                                    |
//| 565+E | 1228 | W0 DATA | TCCl0.12_V_1 te=te:565 scalarw(3) @_SINT/CC/MAPR10NoCE3_ARA0 te=te:565 write(0, 0) |
//| 567   | 1228 | W1 DATA |                                                                                    |
//| 565   | 1229 | R0 DATA |                                                                                    |
//| 565+E | 1229 | W0 DATA | TCCl0.12_V_1 te=te:565 scalarw(3) @_SINT/CC/MAPR10NoCE2_ARA0 te=te:565 write(0, 0) |
//| 568   | 1229 | W1 DATA |                                                                                    |
//| 565   | 1230 | R0 DATA |                                                                                    |
//| 565+E | 1230 | W0 DATA | TCCl0.12_V_1 te=te:565 scalarw(3) @_SINT/CC/MAPR10NoCE1_ARA0 te=te:565 write(0, 0) |
//| 569   | 1230 | W1 DATA |                                                                                    |
//| 565   | 1231 | R0 DATA |                                                                                    |
//| 565+E | 1231 | W0 DATA | TCCl0.12_V_1 te=te:565 scalarw(3) @_SINT/CC/MAPR10NoCE0_ARA0 te=te:565 write(0, 0) |
//| 570   | 1231 | W1 DATA |                                                                                    |
//| 565   | 1232 | R0 DATA |                                                                                    |
//| 565+E | 1232 | W0 DATA | TCCl0.12_V_1 te=te:565 scalarw(4) TCCl0.12_V_0 te=te:565 scalarw(1+TCCl0.12_V_0)   |
//*-------+------+---------+------------------------------------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X109:"xpc10:109" 1237 :  major_start_pcl=571   edge_private_start/end=-1/-1 exec=571 (dend=0)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X109:"xpc10:109" 1236 :  major_start_pcl=571   edge_private_start/end=575/575 exec=571 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X109:"xpc10:109" 1235 :  major_start_pcl=571   edge_private_start/end=574/574 exec=571 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X109:"xpc10:109" 1234 :  major_start_pcl=571   edge_private_start/end=573/573 exec=571 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X109:"xpc10:109" 1233 :  major_start_pcl=571   edge_private_start/end=572/572 exec=571 (dend=1)
//Simple greedy schedule for res2: Thread=xpc10 state=X109:"xpc10:109"
//res2: Thread=xpc10 state=X109:"xpc10:109"
//*-------+------+---------+------------------------------------------------------------------------------------*
//| pc    | eno  | Phaser  | Work                                                                               |
//*-------+------+---------+------------------------------------------------------------------------------------*
//| 571   | -    | R0 CTRL |                                                                                    |
//| 571   | 1233 | R0 DATA |                                                                                    |
//| 571+E | 1233 | W0 DATA | TCCl0.12_V_1 te=te:571 scalarw(3) @_SINT/CC/MAPR10NoCE3_ARA0 te=te:571 write(0, 0) |
//| 572   | 1233 | W1 DATA |                                                                                    |
//| 571   | 1234 | R0 DATA |                                                                                    |
//| 571+E | 1234 | W0 DATA | TCCl0.12_V_1 te=te:571 scalarw(3) @_SINT/CC/MAPR10NoCE2_ARA0 te=te:571 write(0, 0) |
//| 573   | 1234 | W1 DATA |                                                                                    |
//| 571   | 1235 | R0 DATA |                                                                                    |
//| 571+E | 1235 | W0 DATA | TCCl0.12_V_1 te=te:571 scalarw(3) @_SINT/CC/MAPR10NoCE1_ARA0 te=te:571 write(0, 0) |
//| 574   | 1235 | W1 DATA |                                                                                    |
//| 571   | 1236 | R0 DATA |                                                                                    |
//| 571+E | 1236 | W0 DATA | TCCl0.12_V_1 te=te:571 scalarw(3) @_SINT/CC/MAPR10NoCE0_ARA0 te=te:571 write(0, 0) |
//| 575   | 1236 | W1 DATA |                                                                                    |
//| 571   | 1237 | R0 DATA |                                                                                    |
//| 571+E | 1237 | W0 DATA | TCCl0.12_V_1 te=te:571 scalarw(4) TCCl0.12_V_0 te=te:571 scalarw(1+TCCl0.12_V_0)   |
//*-------+------+---------+------------------------------------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X110:"xpc10:110" 1249 :  major_start_pcl=576   edge_private_start/end=-1/-1 exec=576 (dend=0)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X110:"xpc10:110" 1248 :  major_start_pcl=576   edge_private_start/end=587/587 exec=576 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X110:"xpc10:110" 1247 :  major_start_pcl=576   edge_private_start/end=586/586 exec=576 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X110:"xpc10:110" 1246 :  major_start_pcl=576   edge_private_start/end=585/585 exec=576 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X110:"xpc10:110" 1245 :  major_start_pcl=576   edge_private_start/end=584/584 exec=576 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X110:"xpc10:110" 1244 :  major_start_pcl=576   edge_private_start/end=583/583 exec=576 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X110:"xpc10:110" 1243 :  major_start_pcl=576   edge_private_start/end=582/582 exec=576 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X110:"xpc10:110" 1242 :  major_start_pcl=576   edge_private_start/end=581/581 exec=576 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X110:"xpc10:110" 1241 :  major_start_pcl=576   edge_private_start/end=580/580 exec=576 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X110:"xpc10:110" 1240 :  major_start_pcl=576   edge_private_start/end=579/579 exec=576 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X110:"xpc10:110" 1239 :  major_start_pcl=576   edge_private_start/end=578/578 exec=576 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X110:"xpc10:110" 1238 :  major_start_pcl=576   edge_private_start/end=577/577 exec=576 (dend=1)
//Simple greedy schedule for res2: Thread=xpc10 state=X110:"xpc10:110"
//res2: Thread=xpc10 state=X110:"xpc10:110"
//*-------+------+---------+------------------------------------------------------------------------------------*
//| pc    | eno  | Phaser  | Work                                                                               |
//*-------+------+---------+------------------------------------------------------------------------------------*
//| 576   | -    | R0 CTRL |                                                                                    |
//| 576   | 1238 | R0 DATA |                                                                                    |
//| 576+E | 1238 | W0 DATA | TCCl0.12_V_1 te=te:576 scalarw(2) @_SINT/CC/MAPR10NoCE2_ARA0 te=te:576 write(0, 0) |
//| 577   | 1238 | W1 DATA |                                                                                    |
//| 576   | 1239 | R0 DATA |                                                                                    |
//| 576+E | 1239 | W0 DATA | TCCl0.12_V_1 te=te:576 scalarw(2) @_SINT/CC/MAPR10NoCE1_ARA0 te=te:576 write(0, 0) |
//| 578   | 1239 | W1 DATA |                                                                                    |
//| 576   | 1240 | R0 DATA |                                                                                    |
//| 576+E | 1240 | W0 DATA | TCCl0.12_V_1 te=te:576 scalarw(2) @_SINT/CC/MAPR10NoCE0_ARA0 te=te:576 write(0, 0) |
//| 579   | 1240 | W1 DATA |                                                                                    |
//| 576   | 1241 | R0 DATA |                                                                                    |
//| 576+E | 1241 | W0 DATA | TCCl0.12_V_1 te=te:576 scalarw(2) @_SINT/CC/MAPR10NoCE3_ARA0 te=te:576 write(0, 0) |
//| 580   | 1241 | W1 DATA |                                                                                    |
//| 576   | 1242 | R0 DATA |                                                                                    |
//| 576+E | 1242 | W0 DATA | TCCl0.12_V_1 te=te:576 scalarw(2) @_SINT/CC/MAPR10NoCE2_ARA0 te=te:576 write(0, 0) |
//| 581   | 1242 | W1 DATA |                                                                                    |
//| 576   | 1243 | R0 DATA |                                                                                    |
//| 576+E | 1243 | W0 DATA | TCCl0.12_V_1 te=te:576 scalarw(2) @_SINT/CC/MAPR10NoCE1_ARA0 te=te:576 write(0, 0) |
//| 582   | 1243 | W1 DATA |                                                                                    |
//| 576   | 1244 | R0 DATA |                                                                                    |
//| 576+E | 1244 | W0 DATA | TCCl0.12_V_1 te=te:576 scalarw(2) @_SINT/CC/MAPR10NoCE0_ARA0 te=te:576 write(0, 0) |
//| 583   | 1244 | W1 DATA |                                                                                    |
//| 576   | 1245 | R0 DATA |                                                                                    |
//| 576+E | 1245 | W0 DATA | TCCl0.12_V_1 te=te:576 scalarw(3) @_SINT/CC/MAPR10NoCE3_ARA0 te=te:576 write(0, 0) |
//| 584   | 1245 | W1 DATA |                                                                                    |
//| 576   | 1246 | R0 DATA |                                                                                    |
//| 576+E | 1246 | W0 DATA | TCCl0.12_V_1 te=te:576 scalarw(3) @_SINT/CC/MAPR10NoCE2_ARA0 te=te:576 write(0, 0) |
//| 585   | 1246 | W1 DATA |                                                                                    |
//| 576   | 1247 | R0 DATA |                                                                                    |
//| 576+E | 1247 | W0 DATA | TCCl0.12_V_1 te=te:576 scalarw(3) @_SINT/CC/MAPR10NoCE1_ARA0 te=te:576 write(0, 0) |
//| 586   | 1247 | W1 DATA |                                                                                    |
//| 576   | 1248 | R0 DATA |                                                                                    |
//| 576+E | 1248 | W0 DATA | TCCl0.12_V_1 te=te:576 scalarw(3) @_SINT/CC/MAPR10NoCE0_ARA0 te=te:576 write(0, 0) |
//| 587   | 1248 | W1 DATA |                                                                                    |
//| 576   | 1249 | R0 DATA |                                                                                    |
//| 576+E | 1249 | W0 DATA | TCCl0.12_V_1 te=te:576 scalarw(4) TCCl0.12_V_0 te=te:576 scalarw(1+TCCl0.12_V_0)   |
//*-------+------+---------+------------------------------------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X111:"xpc10:111" 1260 :  major_start_pcl=588   edge_private_start/end=-1/-1 exec=588 (dend=0)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X111:"xpc10:111" 1259 :  major_start_pcl=588   edge_private_start/end=598/598 exec=588 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X111:"xpc10:111" 1258 :  major_start_pcl=588   edge_private_start/end=597/597 exec=588 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X111:"xpc10:111" 1257 :  major_start_pcl=588   edge_private_start/end=596/596 exec=588 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X111:"xpc10:111" 1256 :  major_start_pcl=588   edge_private_start/end=595/595 exec=588 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X111:"xpc10:111" 1255 :  major_start_pcl=588   edge_private_start/end=594/594 exec=588 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X111:"xpc10:111" 1254 :  major_start_pcl=588   edge_private_start/end=593/593 exec=588 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X111:"xpc10:111" 1253 :  major_start_pcl=588   edge_private_start/end=592/592 exec=588 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X111:"xpc10:111" 1252 :  major_start_pcl=588   edge_private_start/end=591/591 exec=588 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X111:"xpc10:111" 1251 :  major_start_pcl=588   edge_private_start/end=590/590 exec=588 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X111:"xpc10:111" 1250 :  major_start_pcl=588   edge_private_start/end=589/589 exec=588 (dend=1)
//Simple greedy schedule for res2: Thread=xpc10 state=X111:"xpc10:111"
//res2: Thread=xpc10 state=X111:"xpc10:111"
//*-------+------+---------+------------------------------------------------------------------------------------*
//| pc    | eno  | Phaser  | Work                                                                               |
//*-------+------+---------+------------------------------------------------------------------------------------*
//| 588   | -    | R0 CTRL |                                                                                    |
//| 588   | 1250 | R0 DATA |                                                                                    |
//| 588+E | 1250 | W0 DATA | TCCl0.12_V_1 te=te:588 scalarw(2) @_SINT/CC/MAPR10NoCE1_ARA0 te=te:588 write(0, 0) |
//| 589   | 1250 | W1 DATA |                                                                                    |
//| 588   | 1251 | R0 DATA |                                                                                    |
//| 588+E | 1251 | W0 DATA | TCCl0.12_V_1 te=te:588 scalarw(2) @_SINT/CC/MAPR10NoCE0_ARA0 te=te:588 write(0, 0) |
//| 590   | 1251 | W1 DATA |                                                                                    |
//| 588   | 1252 | R0 DATA |                                                                                    |
//| 588+E | 1252 | W0 DATA | TCCl0.12_V_1 te=te:588 scalarw(2) @_SINT/CC/MAPR10NoCE3_ARA0 te=te:588 write(0, 0) |
//| 591   | 1252 | W1 DATA |                                                                                    |
//| 588   | 1253 | R0 DATA |                                                                                    |
//| 588+E | 1253 | W0 DATA | TCCl0.12_V_1 te=te:588 scalarw(2) @_SINT/CC/MAPR10NoCE2_ARA0 te=te:588 write(0, 0) |
//| 592   | 1253 | W1 DATA |                                                                                    |
//| 588   | 1254 | R0 DATA |                                                                                    |
//| 588+E | 1254 | W0 DATA | TCCl0.12_V_1 te=te:588 scalarw(2) @_SINT/CC/MAPR10NoCE1_ARA0 te=te:588 write(0, 0) |
//| 593   | 1254 | W1 DATA |                                                                                    |
//| 588   | 1255 | R0 DATA |                                                                                    |
//| 588+E | 1255 | W0 DATA | TCCl0.12_V_1 te=te:588 scalarw(2) @_SINT/CC/MAPR10NoCE0_ARA0 te=te:588 write(0, 0) |
//| 594   | 1255 | W1 DATA |                                                                                    |
//| 588   | 1256 | R0 DATA |                                                                                    |
//| 588+E | 1256 | W0 DATA | TCCl0.12_V_1 te=te:588 scalarw(3) @_SINT/CC/MAPR10NoCE3_ARA0 te=te:588 write(0, 0) |
//| 595   | 1256 | W1 DATA |                                                                                    |
//| 588   | 1257 | R0 DATA |                                                                                    |
//| 588+E | 1257 | W0 DATA | TCCl0.12_V_1 te=te:588 scalarw(3) @_SINT/CC/MAPR10NoCE2_ARA0 te=te:588 write(0, 0) |
//| 596   | 1257 | W1 DATA |                                                                                    |
//| 588   | 1258 | R0 DATA |                                                                                    |
//| 588+E | 1258 | W0 DATA | TCCl0.12_V_1 te=te:588 scalarw(3) @_SINT/CC/MAPR10NoCE1_ARA0 te=te:588 write(0, 0) |
//| 597   | 1258 | W1 DATA |                                                                                    |
//| 588   | 1259 | R0 DATA |                                                                                    |
//| 588+E | 1259 | W0 DATA | TCCl0.12_V_1 te=te:588 scalarw(3) @_SINT/CC/MAPR10NoCE0_ARA0 te=te:588 write(0, 0) |
//| 598   | 1259 | W1 DATA |                                                                                    |
//| 588   | 1260 | R0 DATA |                                                                                    |
//| 588+E | 1260 | W0 DATA | TCCl0.12_V_1 te=te:588 scalarw(4) TCCl0.12_V_0 te=te:588 scalarw(1+TCCl0.12_V_0)   |
//*-------+------+---------+------------------------------------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X112:"xpc10:112" 1270 :  major_start_pcl=599   edge_private_start/end=-1/-1 exec=599 (dend=0)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X112:"xpc10:112" 1269 :  major_start_pcl=599   edge_private_start/end=608/608 exec=599 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X112:"xpc10:112" 1268 :  major_start_pcl=599   edge_private_start/end=607/607 exec=599 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X112:"xpc10:112" 1267 :  major_start_pcl=599   edge_private_start/end=606/606 exec=599 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X112:"xpc10:112" 1266 :  major_start_pcl=599   edge_private_start/end=605/605 exec=599 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X112:"xpc10:112" 1265 :  major_start_pcl=599   edge_private_start/end=604/604 exec=599 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X112:"xpc10:112" 1264 :  major_start_pcl=599   edge_private_start/end=603/603 exec=599 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X112:"xpc10:112" 1263 :  major_start_pcl=599   edge_private_start/end=602/602 exec=599 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X112:"xpc10:112" 1262 :  major_start_pcl=599   edge_private_start/end=601/601 exec=599 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X112:"xpc10:112" 1261 :  major_start_pcl=599   edge_private_start/end=600/600 exec=599 (dend=1)
//Simple greedy schedule for res2: Thread=xpc10 state=X112:"xpc10:112"
//res2: Thread=xpc10 state=X112:"xpc10:112"
//*-------+------+---------+------------------------------------------------------------------------------------*
//| pc    | eno  | Phaser  | Work                                                                               |
//*-------+------+---------+------------------------------------------------------------------------------------*
//| 599   | -    | R0 CTRL |                                                                                    |
//| 599   | 1261 | R0 DATA |                                                                                    |
//| 599+E | 1261 | W0 DATA | TCCl0.12_V_1 te=te:599 scalarw(2) @_SINT/CC/MAPR10NoCE0_ARA0 te=te:599 write(0, 0) |
//| 600   | 1261 | W1 DATA |                                                                                    |
//| 599   | 1262 | R0 DATA |                                                                                    |
//| 599+E | 1262 | W0 DATA | TCCl0.12_V_1 te=te:599 scalarw(2) @_SINT/CC/MAPR10NoCE3_ARA0 te=te:599 write(0, 0) |
//| 601   | 1262 | W1 DATA |                                                                                    |
//| 599   | 1263 | R0 DATA |                                                                                    |
//| 599+E | 1263 | W0 DATA | TCCl0.12_V_1 te=te:599 scalarw(2) @_SINT/CC/MAPR10NoCE2_ARA0 te=te:599 write(0, 0) |
//| 602   | 1263 | W1 DATA |                                                                                    |
//| 599   | 1264 | R0 DATA |                                                                                    |
//| 599+E | 1264 | W0 DATA | TCCl0.12_V_1 te=te:599 scalarw(2) @_SINT/CC/MAPR10NoCE1_ARA0 te=te:599 write(0, 0) |
//| 603   | 1264 | W1 DATA |                                                                                    |
//| 599   | 1265 | R0 DATA |                                                                                    |
//| 599+E | 1265 | W0 DATA | TCCl0.12_V_1 te=te:599 scalarw(2) @_SINT/CC/MAPR10NoCE0_ARA0 te=te:599 write(0, 0) |
//| 604   | 1265 | W1 DATA |                                                                                    |
//| 599   | 1266 | R0 DATA |                                                                                    |
//| 599+E | 1266 | W0 DATA | TCCl0.12_V_1 te=te:599 scalarw(3) @_SINT/CC/MAPR10NoCE3_ARA0 te=te:599 write(0, 0) |
//| 605   | 1266 | W1 DATA |                                                                                    |
//| 599   | 1267 | R0 DATA |                                                                                    |
//| 599+E | 1267 | W0 DATA | TCCl0.12_V_1 te=te:599 scalarw(3) @_SINT/CC/MAPR10NoCE2_ARA0 te=te:599 write(0, 0) |
//| 606   | 1267 | W1 DATA |                                                                                    |
//| 599   | 1268 | R0 DATA |                                                                                    |
//| 599+E | 1268 | W0 DATA | TCCl0.12_V_1 te=te:599 scalarw(3) @_SINT/CC/MAPR10NoCE1_ARA0 te=te:599 write(0, 0) |
//| 607   | 1268 | W1 DATA |                                                                                    |
//| 599   | 1269 | R0 DATA |                                                                                    |
//| 599+E | 1269 | W0 DATA | TCCl0.12_V_1 te=te:599 scalarw(3) @_SINT/CC/MAPR10NoCE0_ARA0 te=te:599 write(0, 0) |
//| 608   | 1269 | W1 DATA |                                                                                    |
//| 599   | 1270 | R0 DATA |                                                                                    |
//| 599+E | 1270 | W0 DATA | TCCl0.12_V_1 te=te:599 scalarw(4) TCCl0.12_V_0 te=te:599 scalarw(1+TCCl0.12_V_0)   |
//*-------+------+---------+------------------------------------------------------------------------------------*
//

//----------------------------------------------------------

//Report from restructure2:::
//  Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X113:"xpc10:113" 1279 :  major_start_pcl=609   edge_private_start/end=-1/-1 exec=609 (dend=0)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X113:"xpc10:113" 1278 :  major_start_pcl=609   edge_private_start/end=617/617 exec=609 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X113:"xpc10:113" 1277 :  major_start_pcl=609   edge_private_start/end=616/616 exec=609 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X113:"xpc10:113" 1276 :  major_start_pcl=609   edge_private_start/end=615/615 exec=609 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X113:"xpc10:113" 1275 :  major_start_pcl=609   edge_private_start/end=614/614 exec=609 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X113:"xpc10:113" 1274 :  major_start_pcl=609   edge_private_start/end=613/613 exec=609 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X113:"xpc10:113" 1273 :  major_start_pcl=609   edge_private_start/end=612/612 exec=609 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X113:"xpc10:113" 1272 :  major_start_pcl=609   edge_private_start/end=611/611 exec=609 (dend=1)
//,   Absolute key numbers for scheduled edge res2: Thread=xpc10 state=X113:"xpc10:113" 1271 :  major_start_pcl=609   edge_private_start/end=610/610 exec=609 (dend=1)
//Simple greedy schedule for res2: Thread=xpc10 state=X113:"xpc10:113"
//res2: Thread=xpc10 state=X113:"xpc10:113"
//*-------+------+---------+------------------------------------------------------------------------------------*
//| pc    | eno  | Phaser  | Work                                                                               |
//*-------+------+---------+------------------------------------------------------------------------------------*
//| 609   | -    | R0 CTRL |                                                                                    |
//| 609   | 1271 | R0 DATA |                                                                                    |
//| 609+E | 1271 | W0 DATA | TCCl0.12_V_1 te=te:609 scalarw(2) @_SINT/CC/MAPR10NoCE3_ARA0 te=te:609 write(0, 0) |
//| 610   | 1271 | W1 DATA |                                                                                    |
//| 609   | 1272 | R0 DATA |                                                                                    |
//| 609+E | 1272 | W0 DATA | TCCl0.12_V_1 te=te:609 scalarw(2) @_SINT/CC/MAPR10NoCE2_ARA0 te=te:609 write(0, 0) |
//| 611   | 1272 | W1 DATA |                                                                                    |
//| 609   | 1273 | R0 DATA |                                                                                    |
//| 609+E | 1273 | W0 DATA | TCCl0.12_V_1 te=te:609 scalarw(2) @_SINT/CC/MAPR10NoCE1_ARA0 te=te:609 write(0, 0) |
//| 612   | 1273 | W1 DATA |                                                                                    |
//| 609   | 1274 | R0 DATA |                                                                                    |
//| 609+E | 1274 | W0 DATA | TCCl0.12_V_1 te=te:609 scalarw(2) @_SINT/CC/MAPR10NoCE0_ARA0 te=te:609 write(0, 0) |
//| 613   | 1274 | W1 DATA |                                                                                    |
//| 609   | 1275 | R0 DATA |                                                                                    |
//| 609+E | 1275 | W0 DATA | TCCl0.12_V_1 te=te:609 scalarw(3) @_SINT/CC/MAPR10NoCE3_ARA0 te=te:609 write(0, 0) |
//| 614   | 1275 | W1 DATA |                                                                                    |
//| 609   | 1276 | R0 DATA |                                                                                    |
//| 609+E | 1276 | W0 DATA | TCCl0.12_V_1 te=te:609 scalarw(3) @_SINT/CC/MAPR10NoCE2_ARA0 te=te:609 write(0, 0) |
//| 615   | 1276 | W1 DATA |                                                                                    |
//| 609   | 1277 | R0 DATA |                                                                                    |
//| 609+E | 1277 | W0 DATA | TCCl0.12_V_1 te=te:609 scalarw(3) @_SINT/CC/MAPR10NoCE1_ARA0 te=te:609 write(0, 0) |
//| 616   | 1277 | W1 DATA |                                                                                    |
//| 609   | 1278 | R0 DATA |                                                                                    |
//| 609+E | 1278 | W0 DATA | TCCl0.12_V_1 te=te:609 scalarw(3) @_SINT/CC/MAPR10NoCE0_ARA0 te=te:609 write(0, 0) |
//| 617   | 1278 | W1 DATA |                                                                                    |
//| 609   | 1279 | R0 DATA |                                                                                    |
//| 609+E | 1279 | W0 DATA | TCCl0.12_V_1 te=te:609 scalarw(4) TCCl0.12_V_0 te=te:609 scalarw(1+TCCl0.12_V_0)   |
//*-------+------+---------+------------------------------------------------------------------------------------*
//

//----------------------------------------------------------

//Report from enumbers:::
//Concise expression alias report.
//
//  E1 =.= S32'715136305I+S32'2147001325I*@_SINT/CC/SCALbx28_seed
//
//  E2 =.= C(@_SINT/CC/SCALbx28_seed)
//
//  E3 =.= C64u(@64_US/CC/SCALbx28_dk)
//
//  E4 =.= 1+@_SINT/CC/SCALbx24_stats_lookups
//
//  E5 =.= 1+@_SINT/CC/SCALbx24_stats_lookup_probes
//
//  E6 =.= TTMT4Main_V_11+51*TClo6.9_V_0
//
//  E7 =.= @_SINT/CC/SCALbx24_waycap
//
//  E8 =.= TCha3.10_V_0%@_SINT/CC/SCALbx24_waycap
//
//  E9 =.= C(COND(@$s@_SINT/CC/SCALbx22_ARB0[TClo6.9_V_0]==X3:"MS", @_SINT/CC/MAPR12NoCE3_ARB0[TClo6.9_V_1], COND(@$s@_SINT/CC/SCALbx22_ARB0[TClo6.9_V_0]==X2:"MS", @_SINT/CC/MAPR12NoCE2_ARB0[TClo6.9_V_1], COND(@$s@_SINT/CC/SCALbx22_ARB0[TClo6.9_V_0]==X1:"MS", @_SINT/CC/MAPR12NoCE1_ARB0[TClo6.9_V_1], COND(@$s@_SINT/CC/SCALbx22_ARB0[TClo6.9_V_0]==X0:"MS", @_SINT/CC/MAPR12NoCE0_ARB0[TClo6.9_V_1], *UNDEF)))))
//
//  E10 =.= C64u(@64_US/CC/SCALbx26_ARA0[TClo6.9_V_2])
//
//  E11 =.= C(@_SINT/CC/SCALbx24_next_free)
//
//  E12 =.= 1+@_SINT/CC/SCALbx24_stats_inserts
//
//  E13 =.= 1+@_SINT/CC/SCALbx24_stats_insert_probes
//
//  E14 =.= 1+@_SINT/CC/SCALbx24_stats_insert_evictions
//
//  E15 =.= C(COND(@$s@_SINT/CC/SCALbx20_ARA0[@_SINT/CC/SCALbx24_next_victim]==X3:"MS", @_SINT/CC/MAPR10NoCE3_ARA0[TCin1.9_V_5], COND(@$s@_SINT/CC/SCALbx20_ARA0[@_SINT/CC/SCALbx24_next_victim]==X2:"MS", @_SINT/CC/MAPR10NoCE2_ARA0[TCin1.9_V_5], COND(@$s@_SINT/CC/SCALbx20_ARA0[@_SINT/CC/SCALbx24_next_victim]==X1:"MS", @_SINT/CC/MAPR10NoCE1_ARA0[TCin1.9_V_5], COND(@$s@_SINT/CC/SCALbx20_ARA0[@_SINT/CC/SCALbx24_next_victim]==X0:"MS", @_SINT/CC/MAPR10NoCE0_ARA0[TCin1.9_V_5], *UNDEF)))))
//
//  E16 =.= C(COND(@$s@_SINT/CC/SCALbx22_ARB0[@_SINT/CC/SCALbx24_next_victim]==X3:"MS", @_SINT/CC/MAPR12NoCE3_ARB0[TCin1.9_V_5], COND(@$s@_SINT/CC/SCALbx22_ARB0[@_SINT/CC/SCALbx24_next_victim]==X2:"MS", @_SINT/CC/MAPR12NoCE2_ARB0[TCin1.9_V_5], COND(@$s@_SINT/CC/SCALbx22_ARB0[@_SINT/CC/SCALbx24_next_victim]==X1:"MS", @_SINT/CC/MAPR12NoCE1_ARB0[TCin1.9_V_5], COND(@$s@_SINT/CC/SCALbx22_ARB0[@_SINT/CC/SCALbx24_next_victim]==X0:"MS", @_SINT/CC/MAPR12NoCE0_ARB0[TCin1.9_V_5], *UNDEF)))))
//
//  E17 =.= 1+@_SINT/CC/SCALbx24_next_victim
//
//  E18 =.= TCin1.9_V_0+51*TCin1.9_V_4
//
//  E19 =.= TCha6.10_V_0%@_SINT/CC/SCALbx24_waycap
//
//  E20 =.= @$s@_SINT/CC/SCALbx20_ARA0[0]==X3:"MS"
//
//  E21 =.= @$s@_SINT/CC/SCALbx20_ARA0[0]==X2:"MS"
//
//  E22 =.= @$s@_SINT/CC/SCALbx20_ARA0[0]==X1:"MS"
//
//  E23 =.= @$s@_SINT/CC/SCALbx20_ARA0[0]==X0:"MS"
//
//  E24 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[0]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]==X3:"MS"]}
//
//  E25 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[0]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]==X2:"MS"]}
//
//  E26 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[0]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]==X1:"MS"]}
//
//  E27 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[0]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]==X0:"MS"]}
//
//  E28 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[0]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]==X3:"MS"]}
//
//  E29 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[0]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]==X2:"MS"]}
//
//  E30 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[0]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]==X1:"MS"]}
//
//  E31 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[0]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]==X0:"MS"]}
//
//  E32 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[0]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]==X3:"MS"]}
//
//  E33 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[0]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]==X2:"MS"]}
//
//  E34 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[0]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]==X1:"MS"]}
//
//  E35 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[0]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]==X0:"MS"]}
//
//  E36 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[0]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]!=X0:"MS"]}
//
//  E37 =.= @$s@_SINT/CC/SCALbx20_ARA0[1]==X3:"MS"
//
//  E38 =.= @$s@_SINT/CC/SCALbx20_ARA0[1]==X2:"MS"
//
//  E39 =.= @$s@_SINT/CC/SCALbx20_ARA0[1]==X1:"MS"
//
//  E40 =.= @$s@_SINT/CC/SCALbx20_ARA0[1]==X0:"MS"
//
//  E41 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[1]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]==X3:"MS"]}
//
//  E42 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[1]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]==X2:"MS"]}
//
//  E43 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[1]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]==X1:"MS"]}
//
//  E44 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[1]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]==X0:"MS"]}
//
//  E45 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[1]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]==X3:"MS"]}
//
//  E46 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[1]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]==X2:"MS"]}
//
//  E47 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[1]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]==X1:"MS"]}
//
//  E48 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[1]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]==X0:"MS"]}
//
//  E49 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[1]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]!=X0:"MS"]}
//
//  E50 =.= @$s@_SINT/CC/SCALbx20_ARA0[2]==X3:"MS"
//
//  E51 =.= @$s@_SINT/CC/SCALbx20_ARA0[2]==X2:"MS"
//
//  E52 =.= @$s@_SINT/CC/SCALbx20_ARA0[2]==X1:"MS"
//
//  E53 =.= @$s@_SINT/CC/SCALbx20_ARA0[2]==X0:"MS"
//
//  E54 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[2]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]==X3:"MS"]}
//
//  E55 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[2]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]==X2:"MS"]}
//
//  E56 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[2]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]==X1:"MS"]}
//
//  E57 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[2]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]==X0:"MS"]}
//
//  E58 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[2]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]!=X0:"MS"]}
//
//  E59 =.= @$s@_SINT/CC/SCALbx20_ARA0[3]==X3:"MS"
//
//  E60 =.= @$s@_SINT/CC/SCALbx20_ARA0[3]==X2:"MS"
//
//  E61 =.= @$s@_SINT/CC/SCALbx20_ARA0[3]==X1:"MS"
//
//  E62 =.= @$s@_SINT/CC/SCALbx20_ARA0[3]==X0:"MS"
//
//  E63 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[3]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]!=X0:"MS"]}
//
//  E64 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[0]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]!=X0:"MS", TCCl0.12_V_0<@_SINT/CC/SCALbx24_waycap]}
//
//  E65 =.= TCCl0.12_V_0>=@_SINT/CC/SCALbx24_waycap
//
//  E66 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[0]==X3:"MS", TCCl0.12_V_0<@_SINT/CC/SCALbx24_waycap]}
//
//  E67 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[0]==X2:"MS", TCCl0.12_V_0<@_SINT/CC/SCALbx24_waycap]}
//
//  E68 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[0]==X1:"MS", TCCl0.12_V_0<@_SINT/CC/SCALbx24_waycap]}
//
//  E69 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[0]==X0:"MS", TCCl0.12_V_0<@_SINT/CC/SCALbx24_waycap]}
//
//  E70 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[0]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]==X3:"MS", TCCl0.12_V_0<@_SINT/CC/SCALbx24_waycap]}
//
//  E71 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[0]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]==X2:"MS", TCCl0.12_V_0<@_SINT/CC/SCALbx24_waycap]}
//
//  E72 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[0]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]==X1:"MS", TCCl0.12_V_0<@_SINT/CC/SCALbx24_waycap]}
//
//  E73 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[0]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]==X0:"MS", TCCl0.12_V_0<@_SINT/CC/SCALbx24_waycap]}
//
//  E74 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[0]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]==X3:"MS", TCCl0.12_V_0<@_SINT/CC/SCALbx24_waycap]}
//
//  E75 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[0]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]==X2:"MS", TCCl0.12_V_0<@_SINT/CC/SCALbx24_waycap]}
//
//  E76 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[0]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]==X1:"MS", TCCl0.12_V_0<@_SINT/CC/SCALbx24_waycap]}
//
//  E77 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[0]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]==X0:"MS", TCCl0.12_V_0<@_SINT/CC/SCALbx24_waycap]}
//
//  E78 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[0]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]==X3:"MS", TCCl0.12_V_0<@_SINT/CC/SCALbx24_waycap]}
//
//  E79 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[0]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]==X2:"MS", TCCl0.12_V_0<@_SINT/CC/SCALbx24_waycap]}
//
//  E80 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[0]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]==X1:"MS", TCCl0.12_V_0<@_SINT/CC/SCALbx24_waycap]}
//
//  E81 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[0]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[0]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]==X0:"MS", TCCl0.12_V_0<@_SINT/CC/SCALbx24_waycap]}
//
//  E82 =.= TTMT4Main_V_4>=S32'21845I
//
//  E83 =.= {[TTMT4Main_V_12==TTMT4Main_V_13, !(|-|(C(TCl6._SPILL_256)))]}
//
//  E84 =.= {[TTMT4Main_V_12!=TTMT4Main_V_13, !(|-|(C(TCl6._SPILL_256)))]}
//
//  E85 =.= TTMT4Main_V_10>=S32'21845I
//
//  E86 =.= TTMT4Main_V_10<S32'21845I
//
//  E87 =.= {[|-|isMODULUS10RRh10vld]; [|-|isMODULUS10_rdy]}
//
//  E88 =.= {[TClo6.9_V_0==X4:"US", TTMT4Main_V_11==(COND(@$s@_SINT/CC/SCALbx20_ARA0[TClo6.9_V_0]==X3:"MS", COND(xpc10nz==X237:"US", @_SINT/CC/MAPR10NoCE3_ARA0_RDD0, SINTCCMAPR10NoCE3ARA0RRh10hold), COND(@$s@_SINT/CC/SCALbx20_ARA0[TClo6.9_V_0]==X2:"MS", COND(xpc10nz==X237:"US", @_SINT/CC/MAPR10NoCE2_ARA0_RDD0, SINTCCMAPR10NoCE2ARA0RRh10hold), COND(@$s@_SINT/CC/SCALbx20_ARA0[TClo6.9_V_0]==X1:"MS", COND(xpc10nz==X237:"US", @_SINT/CC/MAPR10NoCE1_ARA0_RDD0, SINTCCMAPR10NoCE1ARA0RRh10hold), COND(@$s@_SINT/CC/SCALbx20_ARA0[TClo6.9_V_0]==X0:"MS", COND(xpc10nz==X237:"US", @_SINT/CC/MAPR10NoCE0_ARA0_RDD0, SINTCCMAPR10NoCE0ARA0RRh10hold), *UNDEF)))))]}
//
//  E89 =.= {[TClo6.9_V_0!=X4:"US", TTMT4Main_V_11==(COND(@$s@_SINT/CC/SCALbx20_ARA0[TClo6.9_V_0]==X3:"MS", COND(xpc10nz==X237:"US", @_SINT/CC/MAPR10NoCE3_ARA0_RDD0, SINTCCMAPR10NoCE3ARA0RRh10hold), COND(@$s@_SINT/CC/SCALbx20_ARA0[TClo6.9_V_0]==X2:"MS", COND(xpc10nz==X237:"US", @_SINT/CC/MAPR10NoCE2_ARA0_RDD0, SINTCCMAPR10NoCE2ARA0RRh10hold), COND(@$s@_SINT/CC/SCALbx20_ARA0[TClo6.9_V_0]==X1:"MS", COND(xpc10nz==X237:"US", @_SINT/CC/MAPR10NoCE1_ARA0_RDD0, SINTCCMAPR10NoCE1ARA0RRh10hold), COND(@$s@_SINT/CC/SCALbx20_ARA0[TClo6.9_V_0]==X0:"MS", COND(xpc10nz==X237:"US", @_SINT/CC/MAPR10NoCE0_ARA0_RDD0, SINTCCMAPR10NoCE0ARA0RRh10hold), *UNDEF)))))]}
//
//  E90 =.= TTMT4Main_V_11!=(COND(@$s@_SINT/CC/SCALbx20_ARA0[TClo6.9_V_0]==X3:"MS", COND(xpc10nz==X237:"US", @_SINT/CC/MAPR10NoCE3_ARA0_RDD0, SINTCCMAPR10NoCE3ARA0RRh10hold), COND(@$s@_SINT/CC/SCALbx20_ARA0[TClo6.9_V_0]==X2:"MS", COND(xpc10nz==X237:"US", @_SINT/CC/MAPR10NoCE2_ARA0_RDD0, SINTCCMAPR10NoCE2ARA0RRh10hold), COND(@$s@_SINT/CC/SCALbx20_ARA0[TClo6.9_V_0]==X1:"MS", COND(xpc10nz==X237:"US", @_SINT/CC/MAPR10NoCE1_ARA0_RDD0, SINTCCMAPR10NoCE1ARA0RRh10hold), COND(@$s@_SINT/CC/SCALbx20_ARA0[TClo6.9_V_0]==X0:"MS", COND(xpc10nz==X237:"US", @_SINT/CC/MAPR10NoCE0_ARA0_RDD0, SINTCCMAPR10NoCE0ARA0RRh10hold), *UNDEF)))))
//
//  E91 =.= {[!(|-|TTMT4Main_V_14), TTMT4Main_V_12==TTMT4Main_V_13]}
//
//  E92 =.= {[!(|-|TTMT4Main_V_14), TTMT4Main_V_12!=TTMT4Main_V_13]}
//
//  E93 =.= {[TClo6.9_V_0>=4, TClo6.9_V_0!=X4:"US"]}
//
//  E94 =.= {[|-|TCin1.9_V_0, @_SINT/CC/SCALbx24_next_free==4*@_SINT/CC/SCALbx24_waycap]}
//
//  E95 =.= {[|-|TCin1.9_V_0, @_SINT/CC/SCALbx24_next_free!=4*@_SINT/CC/SCALbx24_waycap]}
//
//  E96 =.= {[TCin1.9_V_4>=4, TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X3:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]==X3:"MS"]}
//
//  E97 =.= {[TCin1.9_V_4>=4, TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X3:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]==X2:"MS"]}
//
//  E98 =.= {[TCin1.9_V_4>=4, TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X3:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]==X1:"MS"]}
//
//  E99 =.= {[TCin1.9_V_4>=4, TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X3:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]==X0:"MS"]}
//
//  E100 =.= {[TCin1.9_V_4>=4, TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X3:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]!=X3:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]!=X2:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]!=X1:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]!=X0:"MS"]}
//
//  E101 =.= {[TCin1.9_V_4>=4, TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X2:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]==X3:"MS"]}
//
//  E102 =.= {[TCin1.9_V_4>=4, TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X2:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]==X2:"MS"]}
//
//  E103 =.= {[TCin1.9_V_4>=4, TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X2:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]==X1:"MS"]}
//
//  E104 =.= {[TCin1.9_V_4>=4, TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X2:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]==X0:"MS"]}
//
//  E105 =.= {[TCin1.9_V_4>=4, TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X2:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]!=X3:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]!=X2:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]!=X1:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]!=X0:"MS"]}
//
//  E106 =.= {[TCin1.9_V_4>=4, TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X1:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]==X3:"MS"]}
//
//  E107 =.= {[TCin1.9_V_4>=4, TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X1:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]==X2:"MS"]}
//
//  E108 =.= {[TCin1.9_V_4>=4, TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X1:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]==X1:"MS"]}
//
//  E109 =.= {[TCin1.9_V_4>=4, TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X1:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]==X0:"MS"]}
//
//  E110 =.= {[TCin1.9_V_4>=4, TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X1:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]!=X3:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]!=X2:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]!=X1:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]!=X0:"MS"]}
//
//  E111 =.= {[TCin1.9_V_4>=4, TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X0:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]==X3:"MS"]}
//
//  E112 =.= {[TCin1.9_V_4>=4, TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X0:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]==X2:"MS"]}
//
//  E113 =.= {[TCin1.9_V_4>=4, TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X0:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]==X1:"MS"]}
//
//  E114 =.= {[TCin1.9_V_4>=4, TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X0:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]==X0:"MS"]}
//
//  E115 =.= {[TCin1.9_V_4>=4, TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X0:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]!=X3:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]!=X2:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]!=X1:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]!=X0:"MS"]}
//
//  E116 =.= {[TCin1.9_V_4>=4, TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]!=X0:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]==X3:"MS"]}
//
//  E117 =.= {[TCin1.9_V_4>=4, TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]!=X0:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]==X2:"MS"]}
//
//  E118 =.= {[TCin1.9_V_4>=4, TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]!=X0:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]==X1:"MS"]}
//
//  E119 =.= {[TCin1.9_V_4>=4, TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]!=X0:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]==X0:"MS"]}
//
//  E120 =.= {[TCin1.9_V_4>=4, TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]!=X0:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]!=X3:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]!=X2:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]!=X1:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]!=X0:"MS"]}
//
//  E121 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[@_SINT/CC/SCALbx24_next_victim]==X3:"MS", @$s@_SINT/CC/SCALbx22_ARB0[@_SINT/CC/SCALbx24_next_victim]==X3:"MS"]}
//
//  E122 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[@_SINT/CC/SCALbx24_next_victim]==X3:"MS", @$s@_SINT/CC/SCALbx22_ARB0[@_SINT/CC/SCALbx24_next_victim]==X2:"MS"]}
//
//  E123 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[@_SINT/CC/SCALbx24_next_victim]==X3:"MS", @$s@_SINT/CC/SCALbx22_ARB0[@_SINT/CC/SCALbx24_next_victim]==X1:"MS"]}
//
//  E124 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[@_SINT/CC/SCALbx24_next_victim]==X3:"MS", @$s@_SINT/CC/SCALbx22_ARB0[@_SINT/CC/SCALbx24_next_victim]==X0:"MS"]}
//
//  E125 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[@_SINT/CC/SCALbx24_next_victim]==X3:"MS", @$s@_SINT/CC/SCALbx22_ARB0[@_SINT/CC/SCALbx24_next_victim]!=X3:"MS", @$s@_SINT/CC/SCALbx22_ARB0[@_SINT/CC/SCALbx24_next_victim]!=X2:"MS", @$s@_SINT/CC/SCALbx22_ARB0[@_SINT/CC/SCALbx24_next_victim]!=X1:"MS", @$s@_SINT/CC/SCALbx22_ARB0[@_SINT/CC/SCALbx24_next_victim]!=X0:"MS"]}
//
//  E126 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[@_SINT/CC/SCALbx24_next_victim]==X2:"MS", @$s@_SINT/CC/SCALbx22_ARB0[@_SINT/CC/SCALbx24_next_victim]==X3:"MS"]}
//
//  E127 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[@_SINT/CC/SCALbx24_next_victim]==X2:"MS", @$s@_SINT/CC/SCALbx22_ARB0[@_SINT/CC/SCALbx24_next_victim]==X2:"MS"]}
//
//  E128 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[@_SINT/CC/SCALbx24_next_victim]==X2:"MS", @$s@_SINT/CC/SCALbx22_ARB0[@_SINT/CC/SCALbx24_next_victim]==X1:"MS"]}
//
//  E129 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[@_SINT/CC/SCALbx24_next_victim]==X2:"MS", @$s@_SINT/CC/SCALbx22_ARB0[@_SINT/CC/SCALbx24_next_victim]==X0:"MS"]}
//
//  E130 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[@_SINT/CC/SCALbx24_next_victim]==X2:"MS", @$s@_SINT/CC/SCALbx22_ARB0[@_SINT/CC/SCALbx24_next_victim]!=X3:"MS", @$s@_SINT/CC/SCALbx22_ARB0[@_SINT/CC/SCALbx24_next_victim]!=X2:"MS", @$s@_SINT/CC/SCALbx22_ARB0[@_SINT/CC/SCALbx24_next_victim]!=X1:"MS", @$s@_SINT/CC/SCALbx22_ARB0[@_SINT/CC/SCALbx24_next_victim]!=X0:"MS"]}
//
//  E131 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[@_SINT/CC/SCALbx24_next_victim]==X1:"MS", @$s@_SINT/CC/SCALbx22_ARB0[@_SINT/CC/SCALbx24_next_victim]==X3:"MS"]}
//
//  E132 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[@_SINT/CC/SCALbx24_next_victim]==X1:"MS", @$s@_SINT/CC/SCALbx22_ARB0[@_SINT/CC/SCALbx24_next_victim]==X2:"MS"]}
//
//  E133 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[@_SINT/CC/SCALbx24_next_victim]==X1:"MS", @$s@_SINT/CC/SCALbx22_ARB0[@_SINT/CC/SCALbx24_next_victim]==X1:"MS"]}
//
//  E134 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[@_SINT/CC/SCALbx24_next_victim]==X1:"MS", @$s@_SINT/CC/SCALbx22_ARB0[@_SINT/CC/SCALbx24_next_victim]==X0:"MS"]}
//
//  E135 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[@_SINT/CC/SCALbx24_next_victim]==X1:"MS", @$s@_SINT/CC/SCALbx22_ARB0[@_SINT/CC/SCALbx24_next_victim]!=X3:"MS", @$s@_SINT/CC/SCALbx22_ARB0[@_SINT/CC/SCALbx24_next_victim]!=X2:"MS", @$s@_SINT/CC/SCALbx22_ARB0[@_SINT/CC/SCALbx24_next_victim]!=X1:"MS", @$s@_SINT/CC/SCALbx22_ARB0[@_SINT/CC/SCALbx24_next_victim]!=X0:"MS"]}
//
//  E136 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[@_SINT/CC/SCALbx24_next_victim]==X0:"MS", @$s@_SINT/CC/SCALbx22_ARB0[@_SINT/CC/SCALbx24_next_victim]==X3:"MS"]}
//
//  E137 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[@_SINT/CC/SCALbx24_next_victim]==X0:"MS", @$s@_SINT/CC/SCALbx22_ARB0[@_SINT/CC/SCALbx24_next_victim]==X2:"MS"]}
//
//  E138 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[@_SINT/CC/SCALbx24_next_victim]==X0:"MS", @$s@_SINT/CC/SCALbx22_ARB0[@_SINT/CC/SCALbx24_next_victim]==X1:"MS"]}
//
//  E139 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[@_SINT/CC/SCALbx24_next_victim]==X0:"MS", @$s@_SINT/CC/SCALbx22_ARB0[@_SINT/CC/SCALbx24_next_victim]==X0:"MS"]}
//
//  E140 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[@_SINT/CC/SCALbx24_next_victim]==X0:"MS", @$s@_SINT/CC/SCALbx22_ARB0[@_SINT/CC/SCALbx24_next_victim]!=X3:"MS", @$s@_SINT/CC/SCALbx22_ARB0[@_SINT/CC/SCALbx24_next_victim]!=X2:"MS", @$s@_SINT/CC/SCALbx22_ARB0[@_SINT/CC/SCALbx24_next_victim]!=X1:"MS", @$s@_SINT/CC/SCALbx22_ARB0[@_SINT/CC/SCALbx24_next_victim]!=X0:"MS"]}
//
//  E141 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[@_SINT/CC/SCALbx24_next_victim]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[@_SINT/CC/SCALbx24_next_victim]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[@_SINT/CC/SCALbx24_next_victim]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[@_SINT/CC/SCALbx24_next_victim]!=X0:"MS", @$s@_SINT/CC/SCALbx22_ARB0[@_SINT/CC/SCALbx24_next_victim]==X3:"MS"]}
//
//  E142 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[@_SINT/CC/SCALbx24_next_victim]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[@_SINT/CC/SCALbx24_next_victim]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[@_SINT/CC/SCALbx24_next_victim]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[@_SINT/CC/SCALbx24_next_victim]!=X0:"MS", @$s@_SINT/CC/SCALbx22_ARB0[@_SINT/CC/SCALbx24_next_victim]==X2:"MS"]}
//
//  E143 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[@_SINT/CC/SCALbx24_next_victim]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[@_SINT/CC/SCALbx24_next_victim]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[@_SINT/CC/SCALbx24_next_victim]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[@_SINT/CC/SCALbx24_next_victim]!=X0:"MS", @$s@_SINT/CC/SCALbx22_ARB0[@_SINT/CC/SCALbx24_next_victim]==X1:"MS"]}
//
//  E144 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[@_SINT/CC/SCALbx24_next_victim]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[@_SINT/CC/SCALbx24_next_victim]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[@_SINT/CC/SCALbx24_next_victim]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[@_SINT/CC/SCALbx24_next_victim]!=X0:"MS", @$s@_SINT/CC/SCALbx22_ARB0[@_SINT/CC/SCALbx24_next_victim]==X0:"MS"]}
//
//  E145 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[@_SINT/CC/SCALbx24_next_victim]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[@_SINT/CC/SCALbx24_next_victim]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[@_SINT/CC/SCALbx24_next_victim]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[@_SINT/CC/SCALbx24_next_victim]!=X0:"MS", @$s@_SINT/CC/SCALbx22_ARB0[@_SINT/CC/SCALbx24_next_victim]!=X3:"MS", @$s@_SINT/CC/SCALbx22_ARB0[@_SINT/CC/SCALbx24_next_victim]!=X2:"MS", @$s@_SINT/CC/SCALbx22_ARB0[@_SINT/CC/SCALbx24_next_victim]!=X1:"MS", @$s@_SINT/CC/SCALbx22_ARB0[@_SINT/CC/SCALbx24_next_victim]!=X0:"MS"]}
//
//  E146 =.= @$s@_SINT/CC/SCALbx22_ARB0[@_SINT/CC/SCALbx24_next_victim]==X2:"MS"
//
//  E147 =.= @$s@_SINT/CC/SCALbx22_ARB0[@_SINT/CC/SCALbx24_next_victim]==X1:"MS"
//
//  E148 =.= @$s@_SINT/CC/SCALbx22_ARB0[@_SINT/CC/SCALbx24_next_victim]==X0:"MS"
//
//  E149 =.= {[@$s@_SINT/CC/SCALbx22_ARB0[@_SINT/CC/SCALbx24_next_victim]!=X2:"MS", @$s@_SINT/CC/SCALbx22_ARB0[@_SINT/CC/SCALbx24_next_victim]!=X1:"MS", @$s@_SINT/CC/SCALbx22_ARB0[@_SINT/CC/SCALbx24_next_victim]!=X0:"MS"]}
//
//  E150 =.= {[@$s@_SINT/CC/SCALbx22_ARB0[@_SINT/CC/SCALbx24_next_victim]!=X1:"MS", @$s@_SINT/CC/SCALbx22_ARB0[@_SINT/CC/SCALbx24_next_victim]!=X0:"MS"]}
//
//  E151 =.= @$s@_SINT/CC/SCALbx22_ARB0[@_SINT/CC/SCALbx24_next_victim]!=X0:"MS"
//
//  E152 =.= @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]==X2:"MS"
//
//  E153 =.= @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]==X1:"MS"
//
//  E154 =.= @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]==X0:"MS"
//
//  E155 =.= {[@$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]!=X2:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]!=X1:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]!=X0:"MS"]}
//
//  E156 =.= {[@$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]!=X1:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]!=X0:"MS"]}
//
//  E157 =.= @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]!=X0:"MS"
//
//  E158 =.= {[TCin1.9_V_4==X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X3:"MS", xpc10nz==X473:"US", !(|-|@_SINT/CC/MAPR10NoCE3_ARA0_RDD0)]; [TCin1.9_V_4==X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X3:"MS", xpc10nz!=X473:"US", !(|-|SINTCCMAPR10NoCE3ARA0RRh10hold)]}
//
//  E159 =.= {[TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X3:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]==X3:"MS", xpc10nz==X473:"US", !(|-|@_SINT/CC/MAPR10NoCE3_ARA0_RDD0)]; [TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X3:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]==X3:"MS", xpc10nz!=X473:"US", !(|-|SINTCCMAPR10NoCE3ARA0RRh10hold)]}
//
//  E160 =.= {[TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X3:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]==X2:"MS", xpc10nz==X473:"US", !(|-|@_SINT/CC/MAPR10NoCE3_ARA0_RDD0)]; [TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X3:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]==X2:"MS", xpc10nz!=X473:"US", !(|-|SINTCCMAPR10NoCE3ARA0RRh10hold)]}
//
//  E161 =.= {[TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X3:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]==X1:"MS", xpc10nz==X473:"US", !(|-|@_SINT/CC/MAPR10NoCE3_ARA0_RDD0)]; [TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X3:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]==X1:"MS", xpc10nz!=X473:"US", !(|-|SINTCCMAPR10NoCE3ARA0RRh10hold)]}
//
//  E162 =.= {[TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X3:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]==X0:"MS", xpc10nz==X473:"US", !(|-|@_SINT/CC/MAPR10NoCE3_ARA0_RDD0)]; [TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X3:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]==X0:"MS", xpc10nz!=X473:"US", !(|-|SINTCCMAPR10NoCE3ARA0RRh10hold)]}
//
//  E163 =.= {[TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X3:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]!=X3:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]!=X2:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]!=X1:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]!=X0:"MS", xpc10nz==X473:"US", !(|-|@_SINT/CC/MAPR10NoCE3_ARA0_RDD0)]; [TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X3:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]!=X3:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]!=X2:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]!=X1:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]!=X0:"MS", xpc10nz!=X473:"US", !(|-|SINTCCMAPR10NoCE3ARA0RRh10hold)]}
//
//  E164 =.= {[TCin1.9_V_4==X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X2:"MS", xpc10nz==X473:"US", !(|-|@_SINT/CC/MAPR10NoCE2_ARA0_RDD0)]; [TCin1.9_V_4==X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X2:"MS", xpc10nz!=X473:"US", !(|-|SINTCCMAPR10NoCE2ARA0RRh10hold)]}
//
//  E165 =.= {[TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X2:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]==X3:"MS", xpc10nz==X473:"US", !(|-|@_SINT/CC/MAPR10NoCE2_ARA0_RDD0)]; [TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X2:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]==X3:"MS", xpc10nz!=X473:"US", !(|-|SINTCCMAPR10NoCE2ARA0RRh10hold)]}
//
//  E166 =.= {[TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X2:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]==X2:"MS", xpc10nz==X473:"US", !(|-|@_SINT/CC/MAPR10NoCE2_ARA0_RDD0)]; [TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X2:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]==X2:"MS", xpc10nz!=X473:"US", !(|-|SINTCCMAPR10NoCE2ARA0RRh10hold)]}
//
//  E167 =.= {[TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X2:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]==X1:"MS", xpc10nz==X473:"US", !(|-|@_SINT/CC/MAPR10NoCE2_ARA0_RDD0)]; [TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X2:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]==X1:"MS", xpc10nz!=X473:"US", !(|-|SINTCCMAPR10NoCE2ARA0RRh10hold)]}
//
//  E168 =.= {[TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X2:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]==X0:"MS", xpc10nz==X473:"US", !(|-|@_SINT/CC/MAPR10NoCE2_ARA0_RDD0)]; [TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X2:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]==X0:"MS", xpc10nz!=X473:"US", !(|-|SINTCCMAPR10NoCE2ARA0RRh10hold)]}
//
//  E169 =.= {[TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X2:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]!=X3:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]!=X2:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]!=X1:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]!=X0:"MS", xpc10nz==X473:"US", !(|-|@_SINT/CC/MAPR10NoCE2_ARA0_RDD0)]; [TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X2:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]!=X3:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]!=X2:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]!=X1:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]!=X0:"MS", xpc10nz!=X473:"US", !(|-|SINTCCMAPR10NoCE2ARA0RRh10hold)]}
//
//  E170 =.= {[TCin1.9_V_4==X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X1:"MS", xpc10nz==X473:"US", !(|-|@_SINT/CC/MAPR10NoCE1_ARA0_RDD0)]; [TCin1.9_V_4==X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X1:"MS", xpc10nz!=X473:"US", !(|-|SINTCCMAPR10NoCE1ARA0RRh10hold)]}
//
//  E171 =.= {[TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X1:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]==X3:"MS", xpc10nz==X473:"US", !(|-|@_SINT/CC/MAPR10NoCE1_ARA0_RDD0)]; [TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X1:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]==X3:"MS", xpc10nz!=X473:"US", !(|-|SINTCCMAPR10NoCE1ARA0RRh10hold)]}
//
//  E172 =.= {[TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X1:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]==X2:"MS", xpc10nz==X473:"US", !(|-|@_SINT/CC/MAPR10NoCE1_ARA0_RDD0)]; [TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X1:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]==X2:"MS", xpc10nz!=X473:"US", !(|-|SINTCCMAPR10NoCE1ARA0RRh10hold)]}
//
//  E173 =.= {[TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X1:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]==X1:"MS", xpc10nz==X473:"US", !(|-|@_SINT/CC/MAPR10NoCE1_ARA0_RDD0)]; [TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X1:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]==X1:"MS", xpc10nz!=X473:"US", !(|-|SINTCCMAPR10NoCE1ARA0RRh10hold)]}
//
//  E174 =.= {[TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X1:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]==X0:"MS", xpc10nz==X473:"US", !(|-|@_SINT/CC/MAPR10NoCE1_ARA0_RDD0)]; [TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X1:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]==X0:"MS", xpc10nz!=X473:"US", !(|-|SINTCCMAPR10NoCE1ARA0RRh10hold)]}
//
//  E175 =.= {[TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X1:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]!=X3:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]!=X2:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]!=X1:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]!=X0:"MS", xpc10nz==X473:"US", !(|-|@_SINT/CC/MAPR10NoCE1_ARA0_RDD0)]; [TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X1:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]!=X3:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]!=X2:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]!=X1:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]!=X0:"MS", xpc10nz!=X473:"US", !(|-|SINTCCMAPR10NoCE1ARA0RRh10hold)]}
//
//  E176 =.= {[TCin1.9_V_4==X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X0:"MS", xpc10nz==X473:"US", !(|-|@_SINT/CC/MAPR10NoCE0_ARA0_RDD0)]; [TCin1.9_V_4==X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X0:"MS", xpc10nz!=X473:"US", !(|-|SINTCCMAPR10NoCE0ARA0RRh10hold)]}
//
//  E177 =.= {[TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X0:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]==X3:"MS", xpc10nz==X473:"US", !(|-|@_SINT/CC/MAPR10NoCE0_ARA0_RDD0)]; [TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X0:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]==X3:"MS", xpc10nz!=X473:"US", !(|-|SINTCCMAPR10NoCE0ARA0RRh10hold)]}
//
//  E178 =.= {[TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X0:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]==X2:"MS", xpc10nz==X473:"US", !(|-|@_SINT/CC/MAPR10NoCE0_ARA0_RDD0)]; [TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X0:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]==X2:"MS", xpc10nz!=X473:"US", !(|-|SINTCCMAPR10NoCE0ARA0RRh10hold)]}
//
//  E179 =.= {[TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X0:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]==X1:"MS", xpc10nz==X473:"US", !(|-|@_SINT/CC/MAPR10NoCE0_ARA0_RDD0)]; [TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X0:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]==X1:"MS", xpc10nz!=X473:"US", !(|-|SINTCCMAPR10NoCE0ARA0RRh10hold)]}
//
//  E180 =.= {[TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X0:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]==X0:"MS", xpc10nz==X473:"US", !(|-|@_SINT/CC/MAPR10NoCE0_ARA0_RDD0)]; [TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X0:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]==X0:"MS", xpc10nz!=X473:"US", !(|-|SINTCCMAPR10NoCE0ARA0RRh10hold)]}
//
//  E181 =.= {[TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X0:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]!=X3:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]!=X2:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]!=X1:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]!=X0:"MS", xpc10nz==X473:"US", !(|-|@_SINT/CC/MAPR10NoCE0_ARA0_RDD0)]; [TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X0:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]!=X3:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]!=X2:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]!=X1:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]!=X0:"MS", xpc10nz!=X473:"US", !(|-|SINTCCMAPR10NoCE0ARA0RRh10hold)]}
//
//  E182 =.= {[TCin1.9_V_4==X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]!=X0:"MS"]}
//
//  E183 =.= {[TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]!=X0:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]==X3:"MS"]}
//
//  E184 =.= {[TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]!=X0:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]==X2:"MS"]}
//
//  E185 =.= {[TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]!=X0:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]==X1:"MS"]}
//
//  E186 =.= {[TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]!=X0:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]==X0:"MS"]}
//
//  E187 =.= {[TCin1.9_V_4!=X4:"US", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]!=X0:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]!=X3:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]!=X2:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]!=X1:"MS", @$s@_SINT/CC/SCALbx22_ARB0[TCin1.9_V_4]!=X0:"MS"]}
//
//  E188 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X3:"MS", xpc10nz==X473:"US", |-|@_SINT/CC/MAPR10NoCE3_ARA0_RDD0]; [@$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X3:"MS", xpc10nz!=X473:"US", |-|SINTCCMAPR10NoCE3ARA0RRh10hold]; [@$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X1:"MS", xpc10nz==X473:"US", |-|@_SINT/CC/MAPR10NoCE1_ARA0_RDD0]; [@$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X1:"MS", xpc10nz!=X473:"US", |-|SINTCCMAPR10NoCE1ARA0RRh10hold]; [@$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X0:"MS", xpc10nz==X473:"US", |-|@_SINT/CC/MAPR10NoCE0_ARA0_RDD0]; [@$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X0:"MS", xpc10nz!=X473:"US", |-|SINTCCMAPR10NoCE0ARA0RRh10hold]; [@$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X2:"MS", xpc10nz==X473:"US", |-|@_SINT/CC/MAPR10NoCE2_ARA0_RDD0]; [@$s@_SINT/CC/SCALbx20_ARA0[TCin1.9_V_4]==X2:"MS", xpc10nz!=X473:"US", |-|SINTCCMAPR10NoCE2ARA0RRh10hold]}
//
//  E189 =.= @$s@_SINT/CC/SCALbx20_ARA0[TCCl0.12_V_1]==X2:"MS"
//
//  E190 =.= @$s@_SINT/CC/SCALbx20_ARA0[TCCl0.12_V_1]==X1:"MS"
//
//  E191 =.= @$s@_SINT/CC/SCALbx20_ARA0[TCCl0.12_V_1]==X0:"MS"
//
//  E192 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[TCCl0.12_V_1]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[TCCl0.12_V_1]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[TCCl0.12_V_1]!=X0:"MS"]}
//
//  E193 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[TCCl0.12_V_1]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[TCCl0.12_V_1]!=X0:"MS"]}
//
//  E194 =.= @$s@_SINT/CC/SCALbx20_ARA0[TCCl0.12_V_1]!=X0:"MS"
//
//  E195 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[3]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]!=X0:"MS"]}
//
//  E196 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[3]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]!=X0:"MS"]}
//
//  E197 =.= @$s@_SINT/CC/SCALbx20_ARA0[3]!=X0:"MS"
//
//  E198 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[2]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]==X3:"MS"]}
//
//  E199 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[2]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]==X2:"MS"]}
//
//  E200 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[2]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]==X1:"MS"]}
//
//  E201 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[2]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]==X0:"MS"]}
//
//  E202 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[2]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]!=X0:"MS"]}
//
//  E203 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[2]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]==X3:"MS"]}
//
//  E204 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[2]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]==X2:"MS"]}
//
//  E205 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[2]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]==X1:"MS"]}
//
//  E206 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[2]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]==X0:"MS"]}
//
//  E207 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[2]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]!=X0:"MS"]}
//
//  E208 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[2]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]==X3:"MS"]}
//
//  E209 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[2]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]==X2:"MS"]}
//
//  E210 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[2]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]==X1:"MS"]}
//
//  E211 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[2]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]==X0:"MS"]}
//
//  E212 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[2]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]!=X0:"MS"]}
//
//  E213 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[1]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]==X3:"MS"]}
//
//  E214 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[1]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]==X2:"MS"]}
//
//  E215 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[1]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]==X1:"MS"]}
//
//  E216 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[1]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]==X0:"MS"]}
//
//  E217 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[1]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]==X3:"MS"]}
//
//  E218 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[1]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]==X2:"MS"]}
//
//  E219 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[1]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]==X1:"MS"]}
//
//  E220 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[1]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]==X0:"MS"]}
//
//  E221 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[1]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]!=X0:"MS"]}
//
//  E222 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[1]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]==X3:"MS"]}
//
//  E223 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[1]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]==X2:"MS"]}
//
//  E224 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[1]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]==X1:"MS"]}
//
//  E225 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[1]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]==X0:"MS"]}
//
//  E226 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[1]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]==X3:"MS"]}
//
//  E227 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[1]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]==X2:"MS"]}
//
//  E228 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[1]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]==X1:"MS"]}
//
//  E229 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[1]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]==X0:"MS"]}
//
//  E230 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[1]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[1]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]!=X0:"MS"]}
//
//  E231 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[1]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]==X3:"MS"]}
//
//  E232 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[1]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]==X2:"MS"]}
//
//  E233 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[1]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]==X1:"MS"]}
//
//  E234 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[1]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]==X0:"MS"]}
//
//  E235 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[1]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]==X3:"MS"]}
//
//  E236 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[1]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]==X2:"MS"]}
//
//  E237 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[1]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]==X1:"MS"]}
//
//  E238 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[1]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]==X0:"MS"]}
//
//  E239 =.= {[@$s@_SINT/CC/SCALbx20_ARA0[1]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[2]!=X0:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]!=X3:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]!=X2:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]!=X1:"MS", @$s@_SINT/CC/SCALbx20_ARA0[3]!=X0:"MS"]}
//

//----------------------------------------------------------

//Report from verilog_render:::
//1 vectors of width 10
//
//28 vectors of width 32
//
//97 vectors of width 1
//
//10 vectors of width 64
//
//1 vectors of width 15
//
//8 vectors of width 13
//
//8 array locations of width 32
//
//928 bits in scalar variables
//
//Total state bits in module = 2946 bits.
//
//354 continuously assigned (wire/non-state) bits 
//
//Total number of leaf cells = 0
//

//Major Statistics Report:
//Thread .cctor uid=cctor10 has 2 CIL instructions in 1 basic blocks
//Thread .cctor uid=cctor12 has 2 CIL instructions in 1 basic blocks
//Thread .cctor uid=cctor14 has 1 CIL instructions in 1 basic blocks
//Thread Main uid=Main10 has 201 CIL instructions in 52 basic blocks
//Thread mpc10 has 114 bevelab control states (pauses)
//Reindexed thread xpc10 with 618 minor control states
// eof (HPR L/S Verilog)
