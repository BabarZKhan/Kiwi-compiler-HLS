

// CBG Orangepath HPR L/S System

// Verilog output file generated at 21/03/2016 11:19:37
// Kiwi Scientific Acceleration (KiwiC .net/CIL/C# to Verilog/SystemC compiler): Version alpha 2.05: 15-Mar-2016 Unix 3.19.8.100
//  /home/djg11/d320/hprls/kiwipro/kiwic/distro/lib/kiwic.exe -vnl-roundtrip=disable -report-each-step -kiwic-finish=enable -kiwic-kcode-dump=enable -log-dir-name=d_obj_sw_test_b sw_test.exe -vnl=sw_test -vnl-rootmodname=DUT -vnl-resets=synchronous
`timescale 1ns/10ps


module DUT(    output [31:0] result,
    output reg signed [63:0] d_monitor,
    output reg [31:0] phase,
    output hf1_dram0bank_opreq,
    input hf1_dram0bank_oprdy,
    input hf1_dram0bank_ack,
    output hf1_dram0bank_rwbar,
    output [255:0] hf1_dram0bank_wdata,
    output [21:0] hf1_dram0bank_addr,
    input [255:0] hf1_dram0bank_rdata,
    output [31:0] hf1_dram0bank_lanes,
    input clk,
    input reset);
  integer TSPru0_12_V_0;
  integer TSPru0_12_V_1;
  integer TSPin0_6_V_0;
  integer TSPen1_8_V_0;
  integer TSPsw1_2_V_0;
  integer TSPsw1_2_V_1;
  integer TSPne2_10_V_0;
  integer TSPne2_10_V_1;
  integer TSPne2_10_V_2;
  integer TSPne2_10_V_3;
  integer TSPne2_10_V_4;
  reg signed [63:0] TSPne2_10_V_7;
  integer TSPen0_17_V_0;
  integer TSPte2_13_V_0;
  integer TSPte2_13_V_1;
  integer TSPte2_13_V_2;
  integer TSPcr2_16_V_0;
  integer TSPcr2_16_V_1;
  reg signed [63:0] TSPcr2_16_V_2;
  reg [7:0] TCpr0_13_V_0;
  reg [7:0] TCpr0_21_V_0;
  reg [7:0] TCpr0_29_V_0;
  reg [7:0] TCpr0_35_V_0;
  reg [7:0] TCpr0_40_V_0;
  reg [7:0] TCpr0_44_V_0;
  integer TSPe1_SPILL_256;
  integer TSPe0_SPILL_256;
  reg [31:0] A_UINT_CC_SCALbx36_crc_reg;
  reg [31:0] A_UINT_CC_SCALbx36_byteno;
  reg [31:0] A_UINT_CC_SCALbx38_byteno;
  reg [31:0] A_UINT_CC_SCALbx38_crc_reg;
  reg signed [31:0] A_SINT_CC_SCALbx32_d2dim0;
  reg signed [31:0] A_SINT_CC_SCALbx44_d2dim0;
  reg signed [31:0] A_SINT_CC_SCALbx40_d2dim0;
  reg signed [31:0] A_SINT_CC_SCALbx46_d2dim0;
  reg signed [31:0] A_SINT_CC_SCALbx42_d2dim0;
  wire [31:0] A_UINT_CC_SCALbx34_ARA0_RDD0;
  reg [8:0] A_UINT_CC_SCALbx34_ARA0_AD0;
  reg A_UINT_CC_SCALbx34_ARA0_WEN0;
  reg A_UINT_CC_SCALbx34_ARA0_REN0;
  reg [31:0] A_UINT_CC_SCALbx34_ARA0_WRD0;
  wire [31:0] A_SINT_CC_SCALbx16_ARA0_RDD0;
  reg [9:0] A_SINT_CC_SCALbx16_ARA0_AD0;
  reg A_SINT_CC_SCALbx16_ARA0_WEN0;
  reg A_SINT_CC_SCALbx16_ARA0_REN0;
  reg [31:0] A_SINT_CC_SCALbx16_ARA0_WRD0;
  wire [15:0] A_16_SS_CC_SCALbx10_ARA0_RDD0;
  reg [7:0] A_16_SS_CC_SCALbx10_ARA0_AD0;
  reg A_16_SS_CC_SCALbx10_ARA0_WEN0;
  reg A_16_SS_CC_SCALbx10_ARA0_REN0;
  reg [15:0] A_16_SS_CC_SCALbx10_ARA0_WRD0;
  wire [15:0] A_16_SS_CC_SCALbx14_ARC0_RDD0;
  reg [7:0] A_16_SS_CC_SCALbx14_ARC0_AD0;
  reg A_16_SS_CC_SCALbx14_ARC0_WEN0;
  reg A_16_SS_CC_SCALbx14_ARC0_REN0;
  reg [15:0] A_16_SS_CC_SCALbx14_ARC0_WRD0;
  wire [15:0] A_16_SS_CC_SCALbx12_ARB0_RDD0;
  reg [5:0] A_16_SS_CC_SCALbx12_ARB0_AD0;
  reg A_16_SS_CC_SCALbx12_ARB0_WEN0;
  reg A_16_SS_CC_SCALbx12_ARB0_REN0;
  reg [15:0] A_16_SS_CC_SCALbx12_ARB0_WRD0;
  wire [31:0] iuMULTIPLIER10_RR;
  reg [31:0] iuMULTIPLIER10_NN;
  reg [31:0] iuMULTIPLIER10_DD;
  wire iuMULTIPLIER10_err;
  wire [63:0] A_64_SS_CC_SCALbx52_ARA0_RDD0;
  reg [7:0] A_64_SS_CC_SCALbx52_ARA0_AD0;
  reg A_64_SS_CC_SCALbx52_ARA0_WEN0;
  reg A_64_SS_CC_SCALbx52_ARA0_REN0;
  reg [63:0] A_64_SS_CC_SCALbx52_ARA0_WRD0;
  wire [31:0] iuMULTIPLIER12_RR;
  reg [31:0] iuMULTIPLIER12_NN;
  reg [31:0] iuMULTIPLIER12_DD;
  wire iuMULTIPLIER12_err;
  wire [63:0] A_64_SS_CC_SCALbx54_ARB0_RDD0;
  reg [7:0] A_64_SS_CC_SCALbx54_ARB0_AD0;
  reg A_64_SS_CC_SCALbx54_ARB0_WEN0;
  reg A_64_SS_CC_SCALbx54_ARB0_REN0;
  reg [63:0] A_64_SS_CC_SCALbx54_ARB0_WRD0;
  wire [31:0] iuMULTIPLIER14_RR;
  reg [31:0] iuMULTIPLIER14_NN;
  reg [31:0] iuMULTIPLIER14_DD;
  wire iuMULTIPLIER14_err;
  wire [63:0] A_64_SS_CC_SCALbx56_ARC0_RDD0;
  reg [7:0] A_64_SS_CC_SCALbx56_ARC0_AD0;
  reg A_64_SS_CC_SCALbx56_ARC0_WEN0;
  reg A_64_SS_CC_SCALbx56_ARC0_REN0;
  reg [63:0] A_64_SS_CC_SCALbx56_ARC0_WRD0;
  wire [63:0] A_64_SS_CC_SCALbx58_ARD0_RDD0;
  reg [7:0] A_64_SS_CC_SCALbx58_ARD0_AD0;
  reg A_64_SS_CC_SCALbx58_ARD0_WEN0;
  reg A_64_SS_CC_SCALbx58_ARD0_REN0;
  reg [63:0] A_64_SS_CC_SCALbx58_ARD0_WRD0;
  wire [31:0] A_SINT_CC_SCALbx26_ARJ0_RDD0;
  reg [6:0] A_SINT_CC_SCALbx26_ARJ0_AD0;
  reg A_SINT_CC_SCALbx26_ARJ0_WEN0;
  wire A_SINT_CC_SCALbx26_ARJ0_REN0;
  reg [31:0] A_SINT_CC_SCALbx26_ARJ0_WRD0;
  reg xpc10_stall;
  wire xpc10_clear;
  reg [15:0] Z16SSCCSCALbx14ARC0RRh10hold;
  reg Z16SSCCSCALbx14ARC0RRh10shot0;
  reg [31:0] UINTCCSCALbx34ARA0RRh12hold;
  reg UINTCCSCALbx34ARA0RRh12shot0;
  reg [31:0] UINTCCSCALbx34ARA0RRh10hold;
  reg UINTCCSCALbx34ARA0RRh10shot0;
  reg [63:0] Z64SSCCSCALbx52ARA0RRh10hold;
  reg Z64SSCCSCALbx52ARA0RRh10shot0;
  reg [63:0] Z64SSCCSCALbx58ARD0RRh10hold;
  reg Z64SSCCSCALbx58ARD0RRh10shot0;
  reg [63:0] Z64SSCCSCALbx56ARC0RRh10hold;
  reg Z64SSCCSCALbx56ARC0RRh10shot0;
  reg [31:0] SINTCCSCALbx16ARA0RRh10hold;
  reg SINTCCSCALbx16ARA0RRh10shot0;
  reg [63:0] Z64SSCCSCALbx54ARB0RRh10hold;
  reg Z64SSCCSCALbx54ARB0RRh10shot0;
  reg [15:0] Z16SSCCSCALbx12ARB0RRh10hold;
  reg Z16SSCCSCALbx12ARB0RRh10shot0;
  reg [15:0] Z16SSCCSCALbx10ARA0RRh10hold;
  reg Z16SSCCSCALbx10ARA0RRh10shot0;
  reg [31:0] iuMULTIPLIER14RRh12hold;
  reg iuMULTIPLIER14RRh12shot0;
  reg iuMULTIPLIER14RRh12shot1;
  reg [31:0] iuMULTIPLIER14RRh10hold;
  reg iuMULTIPLIER14RRh10shot0;
  reg iuMULTIPLIER14RRh10shot1;
  reg [31:0] iuMULTIPLIER12RRh10hold;
  reg iuMULTIPLIER12RRh10shot0;
  reg iuMULTIPLIER12RRh10shot1;
  reg [31:0] iuMULTIPLIER10RRh10hold;
  reg iuMULTIPLIER10RRh10shot0;
  reg iuMULTIPLIER10RRh10shot1;
  reg [8:0] xpc10nz;
 always   @(* )  begin 
       A_SINT_CC_SCALbx26_ARJ0_AD0 = 0;
       A_SINT_CC_SCALbx26_ARJ0_WRD0 = 0;
       A_64_SS_CC_SCALbx58_ARD0_AD0 = 0;
       A_64_SS_CC_SCALbx58_ARD0_WRD0 = 0;
       A_64_SS_CC_SCALbx56_ARC0_AD0 = 0;
       A_64_SS_CC_SCALbx56_ARC0_WRD0 = 0;
       A_64_SS_CC_SCALbx54_ARB0_AD0 = 0;
       A_64_SS_CC_SCALbx54_ARB0_WRD0 = 0;
       A_64_SS_CC_SCALbx52_ARA0_AD0 = 0;
       A_64_SS_CC_SCALbx52_ARA0_WRD0 = 0;
       iuMULTIPLIER14_NN = 0;
       iuMULTIPLIER14_DD = 0;
       iuMULTIPLIER12_NN = 0;
       iuMULTIPLIER12_DD = 0;
       iuMULTIPLIER10_NN = 0;
       iuMULTIPLIER10_DD = 0;
       A_16_SS_CC_SCALbx12_ARB0_AD0 = 0;
       A_16_SS_CC_SCALbx12_ARB0_WRD0 = 0;
       A_16_SS_CC_SCALbx14_ARC0_AD0 = 0;
       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 0;
       A_16_SS_CC_SCALbx10_ARA0_AD0 = 0;
       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 0;
       A_SINT_CC_SCALbx16_ARA0_AD0 = 0;
       A_SINT_CC_SCALbx16_ARA0_WRD0 = 0;
       A_UINT_CC_SCALbx34_ARA0_AD0 = 0;
       A_UINT_CC_SCALbx34_ARA0_WRD0 = 0;
       A_16_SS_CC_SCALbx12_ARB0_REN0 = 0;
       A_16_SS_CC_SCALbx14_ARC0_REN0 = 0;
       A_SINT_CC_SCALbx26_ARJ0_WEN0 = 0;
       A_UINT_CC_SCALbx34_ARA0_REN0 = 0;
       A_64_SS_CC_SCALbx54_ARB0_REN0 = 0;
       A_64_SS_CC_SCALbx58_ARD0_WEN0 = 0;
       A_64_SS_CC_SCALbx58_ARD0_REN0 = 0;
       A_64_SS_CC_SCALbx52_ARA0_REN0 = 0;
       A_64_SS_CC_SCALbx56_ARC0_WEN0 = 0;
       A_64_SS_CC_SCALbx56_ARC0_REN0 = 0;
       A_64_SS_CC_SCALbx54_ARB0_WEN0 = 0;
       A_SINT_CC_SCALbx16_ARA0_REN0 = 0;
       A_64_SS_CC_SCALbx52_ARA0_WEN0 = 0;
       A_16_SS_CC_SCALbx10_ARA0_REN0 = 0;
       A_SINT_CC_SCALbx16_ARA0_WEN0 = 0;
       A_UINT_CC_SCALbx34_ARA0_WEN0 = 0;
       A_16_SS_CC_SCALbx14_ARC0_WEN0 = 0;
       A_16_SS_CC_SCALbx10_ARA0_WEN0 = 0;
       A_16_SS_CC_SCALbx12_ARB0_WEN0 = 0;
      if (!xpc10_stall)  begin 
               A_16_SS_CC_SCALbx12_ARB0_WEN0 = ((xpc10nz==1'd1/*1:US*/) || (xpc10nz==2'd3/*3:US*/) || (xpc10nz==3'd5/*5:US*/) || (xpc10nz
              ==3'd7/*7:US*/) || (xpc10nz==4'd9/*9:US*/) || (xpc10nz==4'd11/*11:US*/) || (xpc10nz==4'd13/*13:US*/) || (xpc10nz==4'd15
              /*15:US*/) || (xpc10nz==5'd17/*17:US*/) || (xpc10nz==5'd19/*19:US*/) || (xpc10nz==5'd18/*18:US*/) || (xpc10nz==5'd16/*16:US*/) || 
              (xpc10nz==4'd14/*14:US*/) || (xpc10nz==4'd12/*12:US*/) || (xpc10nz==4'd10/*10:US*/) || (xpc10nz==4'd8/*8:US*/) || (xpc10nz
              ==3'd6/*6:US*/) || (xpc10nz==3'd4/*4:US*/) || (xpc10nz==2'd2/*2:US*/) || (xpc10nz==0/*0:US*/)? 1'd1: 1'd0);

               A_16_SS_CC_SCALbx10_ARA0_WEN0 = ((xpc10nz==1'd1/*1:US*/) || (xpc10nz==2'd3/*3:US*/) || (xpc10nz==3'd5/*5:US*/) || (xpc10nz
              ==3'd7/*7:US*/) || (xpc10nz==4'd9/*9:US*/) || (xpc10nz==4'd11/*11:US*/) || (xpc10nz==4'd13/*13:US*/) || (xpc10nz==4'd15
              /*15:US*/) || (xpc10nz==5'd17/*17:US*/) || (xpc10nz==5'd19/*19:US*/) || (xpc10nz==5'd21/*21:US*/) || (xpc10nz==5'd23/*23:US*/) || 
              (xpc10nz==5'd25/*25:US*/) || (xpc10nz==5'd27/*27:US*/) || (xpc10nz==5'd29/*29:US*/) || (xpc10nz==5'd31/*31:US*/) || (xpc10nz
              ==6'd33/*33:US*/) || (xpc10nz==6'd35/*35:US*/) || (xpc10nz==6'd37/*37:US*/) || (xpc10nz==6'd39/*39:US*/) || (xpc10nz==6'd41
              /*41:US*/) || (xpc10nz==6'd43/*43:US*/) || (xpc10nz==6'd45/*45:US*/) || (xpc10nz==6'd47/*47:US*/) || (xpc10nz==6'd49/*49:US*/) || 
              (xpc10nz==6'd51/*51:US*/) || (xpc10nz==6'd53/*53:US*/) || (xpc10nz==6'd55/*55:US*/) || (xpc10nz==6'd57/*57:US*/) || (xpc10nz
              ==6'd59/*59:US*/) || (xpc10nz==6'd61/*61:US*/) || (xpc10nz==6'd63/*63:US*/) || (xpc10nz==7'd65/*65:US*/) || (xpc10nz==7'd67
              /*67:US*/) || (xpc10nz==7'd69/*69:US*/) || (xpc10nz==7'd71/*71:US*/) || (xpc10nz==7'd73/*73:US*/) || (xpc10nz==7'd74/*74:US*/) || 
              (xpc10nz==7'd72/*72:US*/) || (xpc10nz==7'd70/*70:US*/) || (xpc10nz==7'd68/*68:US*/) || (xpc10nz==7'd66/*66:US*/) || (xpc10nz
              ==7'd64/*64:US*/) || (xpc10nz==6'd62/*62:US*/) || (xpc10nz==6'd60/*60:US*/) || (xpc10nz==6'd58/*58:US*/) || (xpc10nz==6'd56
              /*56:US*/) || (xpc10nz==6'd54/*54:US*/) || (xpc10nz==6'd52/*52:US*/) || (xpc10nz==6'd50/*50:US*/) || (xpc10nz==6'd48/*48:US*/) || 
              (xpc10nz==6'd46/*46:US*/) || (xpc10nz==6'd44/*44:US*/) || (xpc10nz==6'd42/*42:US*/) || (xpc10nz==6'd40/*40:US*/) || (xpc10nz
              ==6'd38/*38:US*/) || (xpc10nz==6'd36/*36:US*/) || (xpc10nz==6'd34/*34:US*/) || (xpc10nz==6'd32/*32:US*/) || (xpc10nz==5'd30
              /*30:US*/) || (xpc10nz==5'd28/*28:US*/) || (xpc10nz==5'd26/*26:US*/) || (xpc10nz==5'd24/*24:US*/) || (xpc10nz==5'd22/*22:US*/) || 
              (xpc10nz==5'd20/*20:US*/) || (xpc10nz==5'd18/*18:US*/) || (xpc10nz==5'd16/*16:US*/) || (xpc10nz==4'd14/*14:US*/) || (xpc10nz
              ==4'd12/*12:US*/) || (xpc10nz==4'd10/*10:US*/) || (xpc10nz==4'd8/*8:US*/) || (xpc10nz==3'd6/*6:US*/) || (xpc10nz==3'd4/*4:US*/) || 
              (xpc10nz==2'd2/*2:US*/) || (xpc10nz==0/*0:US*/)? 1'd1: 1'd0);

               A_16_SS_CC_SCALbx14_ARC0_WEN0 = ((xpc10nz==1'd1/*1:US*/) || (xpc10nz==2'd3/*3:US*/) || (xpc10nz==3'd5/*5:US*/) || (xpc10nz
              ==3'd7/*7:US*/) || (xpc10nz==4'd9/*9:US*/) || (xpc10nz==4'd11/*11:US*/) || (xpc10nz==4'd13/*13:US*/) || (xpc10nz==4'd15
              /*15:US*/) || (xpc10nz==5'd17/*17:US*/) || (xpc10nz==5'd19/*19:US*/) || (xpc10nz==5'd21/*21:US*/) || (xpc10nz==5'd23/*23:US*/) || 
              (xpc10nz==5'd25/*25:US*/) || (xpc10nz==5'd27/*27:US*/) || (xpc10nz==5'd29/*29:US*/) || (xpc10nz==5'd31/*31:US*/) || (xpc10nz
              ==6'd33/*33:US*/) || (xpc10nz==6'd35/*35:US*/) || (xpc10nz==6'd37/*37:US*/) || (xpc10nz==6'd39/*39:US*/) || (xpc10nz==6'd41
              /*41:US*/) || (xpc10nz==6'd43/*43:US*/) || (xpc10nz==6'd45/*45:US*/) || (xpc10nz==6'd47/*47:US*/) || (xpc10nz==6'd49/*49:US*/) || 
              (xpc10nz==6'd51/*51:US*/) || (xpc10nz==6'd53/*53:US*/) || (xpc10nz==6'd55/*55:US*/) || (xpc10nz==6'd57/*57:US*/) || (xpc10nz
              ==6'd59/*59:US*/) || (xpc10nz==6'd61/*61:US*/) || (xpc10nz==6'd63/*63:US*/) || (xpc10nz==7'd65/*65:US*/) || (xpc10nz==7'd67
              /*67:US*/) || (xpc10nz==7'd69/*69:US*/) || (xpc10nz==7'd71/*71:US*/) || (xpc10nz==7'd73/*73:US*/) || (xpc10nz==7'd75/*75:US*/) || 
              (xpc10nz==7'd76/*76:US*/) || (xpc10nz==7'd74/*74:US*/) || (xpc10nz==7'd72/*72:US*/) || (xpc10nz==7'd70/*70:US*/) || (xpc10nz
              ==7'd68/*68:US*/) || (xpc10nz==7'd66/*66:US*/) || (xpc10nz==7'd64/*64:US*/) || (xpc10nz==6'd62/*62:US*/) || (xpc10nz==6'd60
              /*60:US*/) || (xpc10nz==6'd58/*58:US*/) || (xpc10nz==6'd56/*56:US*/) || (xpc10nz==6'd54/*54:US*/) || (xpc10nz==6'd52/*52:US*/) || 
              (xpc10nz==6'd50/*50:US*/) || (xpc10nz==6'd48/*48:US*/) || (xpc10nz==6'd46/*46:US*/) || (xpc10nz==6'd44/*44:US*/) || (xpc10nz
              ==6'd42/*42:US*/) || (xpc10nz==6'd40/*40:US*/) || (xpc10nz==6'd38/*38:US*/) || (xpc10nz==6'd36/*36:US*/) || (xpc10nz==6'd34
              /*34:US*/) || (xpc10nz==6'd32/*32:US*/) || (xpc10nz==5'd30/*30:US*/) || (xpc10nz==5'd28/*28:US*/) || (xpc10nz==5'd26/*26:US*/) || 
              (xpc10nz==5'd24/*24:US*/) || (xpc10nz==5'd22/*22:US*/) || (xpc10nz==5'd20/*20:US*/) || (xpc10nz==5'd18/*18:US*/) || (xpc10nz
              ==5'd16/*16:US*/) || (xpc10nz==4'd14/*14:US*/) || (xpc10nz==4'd12/*12:US*/) || (xpc10nz==4'd10/*10:US*/) || (xpc10nz==4'd8
              /*8:US*/) || (xpc10nz==3'd6/*6:US*/) || (xpc10nz==3'd4/*4:US*/) || (xpc10nz==2'd2/*2:US*/) || (xpc10nz==0/*0:US*/)? 1'd1
              : 1'd0);

               A_UINT_CC_SCALbx34_ARA0_WEN0 = ((xpc10nz==1'd1/*1:US*/) || (xpc10nz==2'd3/*3:US*/) || (xpc10nz==3'd5/*5:US*/) || (xpc10nz
              ==3'd7/*7:US*/) || (xpc10nz==4'd9/*9:US*/) || (xpc10nz==4'd11/*11:US*/) || (xpc10nz==4'd13/*13:US*/) || (xpc10nz==4'd15
              /*15:US*/) || (xpc10nz==5'd17/*17:US*/) || (xpc10nz==5'd19/*19:US*/) || (xpc10nz==5'd21/*21:US*/) || (xpc10nz==5'd23/*23:US*/) || 
              (xpc10nz==5'd25/*25:US*/) || (xpc10nz==5'd27/*27:US*/) || (xpc10nz==5'd29/*29:US*/) || (xpc10nz==5'd31/*31:US*/) || (xpc10nz
              ==6'd33/*33:US*/) || (xpc10nz==6'd35/*35:US*/) || (xpc10nz==6'd37/*37:US*/) || (xpc10nz==6'd39/*39:US*/) || (xpc10nz==6'd41
              /*41:US*/) || (xpc10nz==6'd43/*43:US*/) || (xpc10nz==6'd45/*45:US*/) || (xpc10nz==6'd47/*47:US*/) || (xpc10nz==6'd49/*49:US*/) || 
              (xpc10nz==6'd51/*51:US*/) || (xpc10nz==6'd53/*53:US*/) || (xpc10nz==6'd55/*55:US*/) || (xpc10nz==6'd57/*57:US*/) || (xpc10nz
              ==6'd59/*59:US*/) || (xpc10nz==6'd61/*61:US*/) || (xpc10nz==6'd63/*63:US*/) || (xpc10nz==7'd65/*65:US*/) || (xpc10nz==7'd67
              /*67:US*/) || (xpc10nz==7'd69/*69:US*/) || (xpc10nz==7'd71/*71:US*/) || (xpc10nz==7'd73/*73:US*/) || (xpc10nz==7'd75/*75:US*/) || 
              (xpc10nz==7'd77/*77:US*/) || (xpc10nz==7'd79/*79:US*/) || (xpc10nz==7'd81/*81:US*/) || (xpc10nz==7'd83/*83:US*/) || (xpc10nz
              ==7'd85/*85:US*/) || (xpc10nz==7'd87/*87:US*/) || (xpc10nz==7'd89/*89:US*/) || (xpc10nz==7'd91/*91:US*/) || (xpc10nz==7'd93
              /*93:US*/) || (xpc10nz==7'd95/*95:US*/) || (xpc10nz==7'd97/*97:US*/) || (xpc10nz==7'd99/*99:US*/) || (xpc10nz==7'd101/*101:US*/) || 
              (xpc10nz==7'd103/*103:US*/) || (xpc10nz==7'd105/*105:US*/) || (xpc10nz==7'd107/*107:US*/) || (xpc10nz==7'd109/*109:US*/) || 
              (xpc10nz==7'd111/*111:US*/) || (xpc10nz==7'd113/*113:US*/) || (xpc10nz==7'd115/*115:US*/) || (xpc10nz==7'd117/*117:US*/) || 
              (xpc10nz==7'd119/*119:US*/) || (xpc10nz==7'd121/*121:US*/) || (xpc10nz==7'd123/*123:US*/) || (xpc10nz==7'd125/*125:US*/) || 
              (xpc10nz==7'd127/*127:US*/) || (xpc10nz==8'd129/*129:US*/) || (xpc10nz==8'd131/*131:US*/) || (xpc10nz==8'd133/*133:US*/) || 
              (xpc10nz==8'd135/*135:US*/) || (xpc10nz==8'd137/*137:US*/) || (xpc10nz==8'd139/*139:US*/) || (xpc10nz==8'd141/*141:US*/) || 
              (xpc10nz==8'd143/*143:US*/) || (xpc10nz==8'd145/*145:US*/) || (xpc10nz==8'd147/*147:US*/) || (xpc10nz==8'd149/*149:US*/) || 
              (xpc10nz==8'd151/*151:US*/) || (xpc10nz==8'd153/*153:US*/) || (xpc10nz==8'd155/*155:US*/) || (xpc10nz==8'd157/*157:US*/) || 
              (xpc10nz==8'd159/*159:US*/) || (xpc10nz==8'd161/*161:US*/) || (xpc10nz==8'd163/*163:US*/) || (xpc10nz==8'd165/*165:US*/) || 
              (xpc10nz==8'd167/*167:US*/) || (xpc10nz==8'd169/*169:US*/) || (xpc10nz==8'd171/*171:US*/) || (xpc10nz==8'd173/*173:US*/) || 
              (xpc10nz==8'd175/*175:US*/) || (xpc10nz==8'd177/*177:US*/) || (xpc10nz==8'd179/*179:US*/) || (xpc10nz==8'd181/*181:US*/) || 
              (xpc10nz==8'd183/*183:US*/) || (xpc10nz==8'd185/*185:US*/) || (xpc10nz==8'd187/*187:US*/) || (xpc10nz==8'd189/*189:US*/) || 
              (xpc10nz==8'd191/*191:US*/) || (xpc10nz==8'd193/*193:US*/) || (xpc10nz==8'd195/*195:US*/) || (xpc10nz==8'd197/*197:US*/) || 
              (xpc10nz==8'd199/*199:US*/) || (xpc10nz==8'd201/*201:US*/) || (xpc10nz==8'd203/*203:US*/) || (xpc10nz==8'd205/*205:US*/) || 
              (xpc10nz==8'd207/*207:US*/) || (xpc10nz==8'd209/*209:US*/) || (xpc10nz==8'd211/*211:US*/) || (xpc10nz==8'd213/*213:US*/) || 
              (xpc10nz==8'd215/*215:US*/) || (xpc10nz==8'd217/*217:US*/) || (xpc10nz==8'd219/*219:US*/) || (xpc10nz==8'd221/*221:US*/) || 
              (xpc10nz==8'd223/*223:US*/) || (xpc10nz==8'd225/*225:US*/) || (xpc10nz==8'd227/*227:US*/) || (xpc10nz==8'd229/*229:US*/) || 
              (xpc10nz==8'd231/*231:US*/) || (xpc10nz==8'd233/*233:US*/) || (xpc10nz==8'd235/*235:US*/) || (xpc10nz==8'd237/*237:US*/) || 
              (xpc10nz==8'd239/*239:US*/) || (xpc10nz==8'd241/*241:US*/) || (xpc10nz==8'd243/*243:US*/) || (xpc10nz==8'd245/*245:US*/) || 
              (xpc10nz==8'd247/*247:US*/) || (xpc10nz==8'd249/*249:US*/) || (xpc10nz==8'd251/*251:US*/) || (xpc10nz==8'd253/*253:US*/) || 
              (xpc10nz==8'd255/*255:US*/) || (xpc10nz==8'd254/*254:US*/) || (xpc10nz==8'd252/*252:US*/) || (xpc10nz==8'd250/*250:US*/) || 
              (xpc10nz==8'd248/*248:US*/) || (xpc10nz==8'd246/*246:US*/) || (xpc10nz==8'd244/*244:US*/) || (xpc10nz==8'd242/*242:US*/) || 
              (xpc10nz==8'd240/*240:US*/) || (xpc10nz==8'd238/*238:US*/) || (xpc10nz==8'd236/*236:US*/) || (xpc10nz==8'd234/*234:US*/) || 
              (xpc10nz==8'd232/*232:US*/) || (xpc10nz==8'd230/*230:US*/) || (xpc10nz==8'd228/*228:US*/) || (xpc10nz==8'd226/*226:US*/) || 
              (xpc10nz==8'd224/*224:US*/) || (xpc10nz==8'd222/*222:US*/) || (xpc10nz==8'd220/*220:US*/) || (xpc10nz==8'd218/*218:US*/) || 
              (xpc10nz==8'd216/*216:US*/) || (xpc10nz==8'd214/*214:US*/) || (xpc10nz==8'd212/*212:US*/) || (xpc10nz==8'd210/*210:US*/) || 
              (xpc10nz==8'd208/*208:US*/) || (xpc10nz==8'd206/*206:US*/) || (xpc10nz==8'd204/*204:US*/) || (xpc10nz==8'd202/*202:US*/) || 
              (xpc10nz==8'd200/*200:US*/) || (xpc10nz==8'd198/*198:US*/) || (xpc10nz==8'd196/*196:US*/) || (xpc10nz==8'd194/*194:US*/) || 
              (xpc10nz==8'd192/*192:US*/) || (xpc10nz==8'd190/*190:US*/) || (xpc10nz==8'd188/*188:US*/) || (xpc10nz==8'd186/*186:US*/) || 
              (xpc10nz==8'd184/*184:US*/) || (xpc10nz==8'd182/*182:US*/) || (xpc10nz==8'd180/*180:US*/) || (xpc10nz==8'd178/*178:US*/) || 
              (xpc10nz==8'd176/*176:US*/) || (xpc10nz==8'd174/*174:US*/) || (xpc10nz==8'd172/*172:US*/) || (xpc10nz==8'd170/*170:US*/) || 
              (xpc10nz==8'd168/*168:US*/) || (xpc10nz==8'd166/*166:US*/) || (xpc10nz==8'd164/*164:US*/) || (xpc10nz==8'd162/*162:US*/) || 
              (xpc10nz==8'd160/*160:US*/) || (xpc10nz==8'd158/*158:US*/) || (xpc10nz==8'd156/*156:US*/) || (xpc10nz==8'd154/*154:US*/) || 
              (xpc10nz==8'd152/*152:US*/) || (xpc10nz==8'd150/*150:US*/) || (xpc10nz==8'd148/*148:US*/) || (xpc10nz==8'd146/*146:US*/) || 
              (xpc10nz==8'd144/*144:US*/) || (xpc10nz==8'd142/*142:US*/) || (xpc10nz==8'd140/*140:US*/) || (xpc10nz==8'd138/*138:US*/) || 
              (xpc10nz==8'd136/*136:US*/) || (xpc10nz==8'd134/*134:US*/) || (xpc10nz==8'd132/*132:US*/) || (xpc10nz==8'd130/*130:US*/) || 
              (xpc10nz==8'd128/*128:US*/) || (xpc10nz==7'd126/*126:US*/) || (xpc10nz==7'd124/*124:US*/) || (xpc10nz==7'd122/*122:US*/) || 
              (xpc10nz==7'd120/*120:US*/) || (xpc10nz==7'd118/*118:US*/) || (xpc10nz==7'd116/*116:US*/) || (xpc10nz==7'd114/*114:US*/) || 
              (xpc10nz==7'd112/*112:US*/) || (xpc10nz==7'd110/*110:US*/) || (xpc10nz==7'd108/*108:US*/) || (xpc10nz==7'd106/*106:US*/) || 
              (xpc10nz==7'd104/*104:US*/) || (xpc10nz==7'd102/*102:US*/) || (xpc10nz==7'd100/*100:US*/) || (xpc10nz==7'd98/*98:US*/) || 
              (xpc10nz==7'd96/*96:US*/) || (xpc10nz==7'd94/*94:US*/) || (xpc10nz==7'd92/*92:US*/) || (xpc10nz==7'd90/*90:US*/) || (xpc10nz
              ==7'd88/*88:US*/) || (xpc10nz==7'd86/*86:US*/) || (xpc10nz==7'd84/*84:US*/) || (xpc10nz==7'd82/*82:US*/) || (xpc10nz==7'd80
              /*80:US*/) || (xpc10nz==7'd78/*78:US*/) || (xpc10nz==7'd76/*76:US*/) || (xpc10nz==7'd74/*74:US*/) || (xpc10nz==7'd72/*72:US*/) || 
              (xpc10nz==7'd70/*70:US*/) || (xpc10nz==7'd68/*68:US*/) || (xpc10nz==7'd66/*66:US*/) || (xpc10nz==7'd64/*64:US*/) || (xpc10nz
              ==6'd62/*62:US*/) || (xpc10nz==6'd60/*60:US*/) || (xpc10nz==6'd58/*58:US*/) || (xpc10nz==6'd56/*56:US*/) || (xpc10nz==6'd54
              /*54:US*/) || (xpc10nz==6'd52/*52:US*/) || (xpc10nz==6'd50/*50:US*/) || (xpc10nz==6'd48/*48:US*/) || (xpc10nz==6'd46/*46:US*/) || 
              (xpc10nz==6'd44/*44:US*/) || (xpc10nz==6'd42/*42:US*/) || (xpc10nz==6'd40/*40:US*/) || (xpc10nz==6'd38/*38:US*/) || (xpc10nz
              ==6'd36/*36:US*/) || (xpc10nz==6'd34/*34:US*/) || (xpc10nz==6'd32/*32:US*/) || (xpc10nz==5'd30/*30:US*/) || (xpc10nz==5'd28
              /*28:US*/) || (xpc10nz==5'd26/*26:US*/) || (xpc10nz==5'd24/*24:US*/) || (xpc10nz==5'd22/*22:US*/) || (xpc10nz==5'd20/*20:US*/) || 
              (xpc10nz==5'd18/*18:US*/) || (xpc10nz==5'd16/*16:US*/) || (xpc10nz==4'd14/*14:US*/) || (xpc10nz==4'd12/*12:US*/) || (xpc10nz
              ==4'd10/*10:US*/) || (xpc10nz==4'd8/*8:US*/) || (xpc10nz==3'd6/*6:US*/) || (xpc10nz==3'd4/*4:US*/) || (xpc10nz==2'd2/*2:US*/) || 
              (xpc10nz==0/*0:US*/)? 1'd1: 1'd0);

               A_SINT_CC_SCALbx16_ARA0_WEN0 = ((xpc10nz==1'd1/*1:US*/) || (xpc10nz==2'd3/*3:US*/) || (xpc10nz==3'd5/*5:US*/) || (xpc10nz
              ==3'd7/*7:US*/) || (xpc10nz==4'd9/*9:US*/) || (xpc10nz==4'd11/*11:US*/) || (xpc10nz==4'd13/*13:US*/) || (xpc10nz==4'd15
              /*15:US*/) || (xpc10nz==5'd17/*17:US*/) || (xpc10nz==5'd19/*19:US*/) || (xpc10nz==5'd21/*21:US*/) || (xpc10nz==5'd23/*23:US*/) || 
              (xpc10nz==5'd25/*25:US*/) || (xpc10nz==5'd27/*27:US*/) || (xpc10nz==5'd29/*29:US*/) || (xpc10nz==5'd31/*31:US*/) || (xpc10nz
              ==6'd33/*33:US*/) || (xpc10nz==6'd35/*35:US*/) || (xpc10nz==6'd37/*37:US*/) || (xpc10nz==6'd39/*39:US*/) || (xpc10nz==6'd41
              /*41:US*/) || (xpc10nz==6'd43/*43:US*/) || (xpc10nz==6'd45/*45:US*/) || (xpc10nz==6'd47/*47:US*/) || (xpc10nz==6'd49/*49:US*/) || 
              (xpc10nz==6'd51/*51:US*/) || (xpc10nz==6'd53/*53:US*/) || (xpc10nz==6'd55/*55:US*/) || (xpc10nz==6'd57/*57:US*/) || (xpc10nz
              ==6'd59/*59:US*/) || (xpc10nz==6'd61/*61:US*/) || (xpc10nz==6'd63/*63:US*/) || (xpc10nz==7'd65/*65:US*/) || (xpc10nz==7'd67
              /*67:US*/) || (xpc10nz==7'd69/*69:US*/) || (xpc10nz==7'd71/*71:US*/) || (xpc10nz==7'd73/*73:US*/) || (xpc10nz==7'd75/*75:US*/) || 
              (xpc10nz==7'd77/*77:US*/) || (xpc10nz==7'd79/*79:US*/) || (xpc10nz==7'd81/*81:US*/) || (xpc10nz==7'd83/*83:US*/) || (xpc10nz
              ==7'd85/*85:US*/) || (xpc10nz==7'd87/*87:US*/) || (xpc10nz==7'd89/*89:US*/) || (xpc10nz==7'd91/*91:US*/) || (xpc10nz==7'd93
              /*93:US*/) || (xpc10nz==7'd95/*95:US*/) || (xpc10nz==7'd97/*97:US*/) || (xpc10nz==7'd99/*99:US*/) || (xpc10nz==7'd101/*101:US*/) || 
              (xpc10nz==7'd103/*103:US*/) || (xpc10nz==7'd105/*105:US*/) || (xpc10nz==7'd107/*107:US*/) || (xpc10nz==7'd109/*109:US*/) || 
              (xpc10nz==7'd111/*111:US*/) || (xpc10nz==7'd113/*113:US*/) || (xpc10nz==7'd115/*115:US*/) || (xpc10nz==7'd117/*117:US*/) || 
              (xpc10nz==7'd119/*119:US*/) || (xpc10nz==7'd121/*121:US*/) || (xpc10nz==7'd123/*123:US*/) || (xpc10nz==7'd125/*125:US*/) || 
              (xpc10nz==7'd127/*127:US*/) || (xpc10nz==8'd129/*129:US*/) || (xpc10nz==8'd131/*131:US*/) || (xpc10nz==8'd133/*133:US*/) || 
              (xpc10nz==8'd135/*135:US*/) || (xpc10nz==8'd137/*137:US*/) || (xpc10nz==8'd139/*139:US*/) || (xpc10nz==8'd141/*141:US*/) || 
              (xpc10nz==8'd143/*143:US*/) || (xpc10nz==8'd145/*145:US*/) || (xpc10nz==8'd147/*147:US*/) || (xpc10nz==8'd149/*149:US*/) || 
              (xpc10nz==8'd151/*151:US*/) || (xpc10nz==8'd153/*153:US*/) || (xpc10nz==8'd155/*155:US*/) || (xpc10nz==8'd157/*157:US*/) || 
              (xpc10nz==8'd159/*159:US*/) || (xpc10nz==8'd161/*161:US*/) || (xpc10nz==8'd163/*163:US*/) || (xpc10nz==8'd165/*165:US*/) || 
              (xpc10nz==8'd167/*167:US*/) || (xpc10nz==8'd169/*169:US*/) || (xpc10nz==8'd171/*171:US*/) || (xpc10nz==8'd173/*173:US*/) || 
              (xpc10nz==8'd175/*175:US*/) || (xpc10nz==8'd177/*177:US*/) || (xpc10nz==8'd179/*179:US*/) || (xpc10nz==8'd181/*181:US*/) || 
              (xpc10nz==8'd183/*183:US*/) || (xpc10nz==8'd185/*185:US*/) || (xpc10nz==8'd187/*187:US*/) || (xpc10nz==8'd189/*189:US*/) || 
              (xpc10nz==8'd191/*191:US*/) || (xpc10nz==8'd193/*193:US*/) || (xpc10nz==8'd195/*195:US*/) || (xpc10nz==8'd197/*197:US*/) || 
              (xpc10nz==8'd199/*199:US*/) || (xpc10nz==8'd201/*201:US*/) || (xpc10nz==8'd203/*203:US*/) || (xpc10nz==8'd205/*205:US*/) || 
              (xpc10nz==8'd207/*207:US*/) || (xpc10nz==8'd209/*209:US*/) || (xpc10nz==8'd211/*211:US*/) || (xpc10nz==8'd213/*213:US*/) || 
              (xpc10nz==8'd215/*215:US*/) || (xpc10nz==8'd217/*217:US*/) || (xpc10nz==8'd219/*219:US*/) || (xpc10nz==8'd221/*221:US*/) || 
              (xpc10nz==8'd223/*223:US*/) || (xpc10nz==8'd225/*225:US*/) || (xpc10nz==8'd227/*227:US*/) || (xpc10nz==8'd229/*229:US*/) || 
              (xpc10nz==8'd231/*231:US*/) || (xpc10nz==8'd233/*233:US*/) || (xpc10nz==8'd235/*235:US*/) || (xpc10nz==8'd237/*237:US*/) || 
              (xpc10nz==8'd239/*239:US*/) || (xpc10nz==8'd241/*241:US*/) || (xpc10nz==8'd243/*243:US*/) || (xpc10nz==8'd245/*245:US*/) || 
              (xpc10nz==8'd247/*247:US*/) || (xpc10nz==8'd249/*249:US*/) || (xpc10nz==8'd251/*251:US*/) || (xpc10nz==8'd253/*253:US*/) || 
              (xpc10nz==8'd255/*255:US*/) || (xpc10nz==9'd257/*257:US*/) || (xpc10nz==9'd259/*259:US*/) || (xpc10nz==9'd261/*261:US*/) || 
              (xpc10nz==9'd263/*263:US*/) || (xpc10nz==9'd265/*265:US*/) || (xpc10nz==9'd267/*267:US*/) || (xpc10nz==9'd269/*269:US*/) || 
              (xpc10nz==9'd271/*271:US*/) || (xpc10nz==9'd273/*273:US*/) || (xpc10nz==9'd275/*275:US*/) || (xpc10nz==9'd277/*277:US*/) || 
              (xpc10nz==9'd279/*279:US*/) || (xpc10nz==9'd281/*281:US*/) || (xpc10nz==9'd283/*283:US*/) || (xpc10nz==9'd285/*285:US*/) || 
              (xpc10nz==9'd287/*287:US*/) || (xpc10nz==9'd289/*289:US*/) || (xpc10nz==9'd291/*291:US*/) || (xpc10nz==9'd293/*293:US*/) || 
              (xpc10nz==9'd295/*295:US*/) || (xpc10nz==9'd297/*297:US*/) || (xpc10nz==9'd299/*299:US*/) || (xpc10nz==9'd301/*301:US*/) || 
              (xpc10nz==9'd303/*303:US*/) || (xpc10nz==9'd305/*305:US*/) || (xpc10nz==9'd307/*307:US*/) || (xpc10nz==9'd309/*309:US*/) || 
              (xpc10nz==9'd311/*311:US*/) || (xpc10nz==9'd313/*313:US*/) || (xpc10nz==9'd315/*315:US*/) || (xpc10nz==9'd317/*317:US*/) || 
              (xpc10nz==9'd319/*319:US*/) || (xpc10nz==9'd321/*321:US*/) || (xpc10nz==9'd323/*323:US*/) || (xpc10nz==9'd325/*325:US*/) || 
              (xpc10nz==9'd327/*327:US*/) || (xpc10nz==9'd329/*329:US*/) || (xpc10nz==9'd331/*331:US*/) || (xpc10nz==9'd333/*333:US*/) || 
              (xpc10nz==9'd335/*335:US*/) || (xpc10nz==9'd337/*337:US*/) || (xpc10nz==9'd339/*339:US*/) || (xpc10nz==9'd341/*341:US*/) || 
              (xpc10nz==9'd343/*343:US*/) || (xpc10nz==9'd345/*345:US*/) || (xpc10nz==9'd347/*347:US*/) || (xpc10nz==9'd349/*349:US*/) || 
              (xpc10nz==9'd351/*351:US*/) || (xpc10nz==9'd353/*353:US*/) || (xpc10nz==9'd355/*355:US*/) || (xpc10nz==9'd357/*357:US*/) || 
              (xpc10nz==9'd359/*359:US*/) || (xpc10nz==9'd361/*361:US*/) || (xpc10nz==9'd363/*363:US*/) || (xpc10nz==9'd365/*365:US*/) || 
              (xpc10nz==9'd367/*367:US*/) || (xpc10nz==9'd369/*369:US*/) || (xpc10nz==9'd371/*371:US*/) || (xpc10nz==9'd373/*373:US*/) || 
              (xpc10nz==9'd375/*375:US*/) || (xpc10nz==9'd377/*377:US*/) || (xpc10nz==9'd379/*379:US*/) || (xpc10nz==9'd381/*381:US*/) || 
              (xpc10nz==9'd383/*383:US*/) || (xpc10nz==9'd385/*385:US*/) || (xpc10nz==9'd387/*387:US*/) || (xpc10nz==9'd389/*389:US*/) || 
              (xpc10nz==9'd391/*391:US*/) || (xpc10nz==9'd393/*393:US*/) || (xpc10nz==9'd395/*395:US*/) || (xpc10nz==9'd397/*397:US*/) || 
              (xpc10nz==9'd399/*399:US*/) || (xpc10nz==9'd398/*398:US*/) || (xpc10nz==9'd396/*396:US*/) || (xpc10nz==9'd394/*394:US*/) || 
              (xpc10nz==9'd392/*392:US*/) || (xpc10nz==9'd390/*390:US*/) || (xpc10nz==9'd388/*388:US*/) || (xpc10nz==9'd386/*386:US*/) || 
              (xpc10nz==9'd384/*384:US*/) || (xpc10nz==9'd382/*382:US*/) || (xpc10nz==9'd380/*380:US*/) || (xpc10nz==9'd378/*378:US*/) || 
              (xpc10nz==9'd376/*376:US*/) || (xpc10nz==9'd374/*374:US*/) || (xpc10nz==9'd372/*372:US*/) || (xpc10nz==9'd370/*370:US*/) || 
              (xpc10nz==9'd368/*368:US*/) || (xpc10nz==9'd366/*366:US*/) || (xpc10nz==9'd364/*364:US*/) || (xpc10nz==9'd362/*362:US*/) || 
              (xpc10nz==9'd360/*360:US*/) || (xpc10nz==9'd358/*358:US*/) || (xpc10nz==9'd356/*356:US*/) || (xpc10nz==9'd354/*354:US*/) || 
              (xpc10nz==9'd352/*352:US*/) || (xpc10nz==9'd350/*350:US*/) || (xpc10nz==9'd348/*348:US*/) || (xpc10nz==9'd346/*346:US*/) || 
              (xpc10nz==9'd344/*344:US*/) || (xpc10nz==9'd342/*342:US*/) || (xpc10nz==9'd340/*340:US*/) || (xpc10nz==9'd338/*338:US*/) || 
              (xpc10nz==9'd336/*336:US*/) || (xpc10nz==9'd334/*334:US*/) || (xpc10nz==9'd332/*332:US*/) || (xpc10nz==9'd330/*330:US*/) || 
              (xpc10nz==9'd328/*328:US*/) || (xpc10nz==9'd326/*326:US*/) || (xpc10nz==9'd324/*324:US*/) || (xpc10nz==9'd322/*322:US*/) || 
              (xpc10nz==9'd320/*320:US*/) || (xpc10nz==9'd318/*318:US*/) || (xpc10nz==9'd316/*316:US*/) || (xpc10nz==9'd314/*314:US*/) || 
              (xpc10nz==9'd312/*312:US*/) || (xpc10nz==9'd310/*310:US*/) || (xpc10nz==9'd308/*308:US*/) || (xpc10nz==9'd306/*306:US*/) || 
              (xpc10nz==9'd304/*304:US*/) || (xpc10nz==9'd302/*302:US*/) || (xpc10nz==9'd300/*300:US*/) || (xpc10nz==9'd298/*298:US*/) || 
              (xpc10nz==9'd296/*296:US*/) || (xpc10nz==9'd294/*294:US*/) || (xpc10nz==9'd292/*292:US*/) || (xpc10nz==9'd290/*290:US*/) || 
              (xpc10nz==9'd288/*288:US*/) || (xpc10nz==9'd286/*286:US*/) || (xpc10nz==9'd284/*284:US*/) || (xpc10nz==9'd282/*282:US*/) || 
              (xpc10nz==9'd280/*280:US*/) || (xpc10nz==9'd278/*278:US*/) || (xpc10nz==9'd276/*276:US*/) || (xpc10nz==9'd274/*274:US*/) || 
              (xpc10nz==9'd272/*272:US*/) || (xpc10nz==9'd270/*270:US*/) || (xpc10nz==9'd268/*268:US*/) || (xpc10nz==9'd266/*266:US*/) || 
              (xpc10nz==9'd264/*264:US*/) || (xpc10nz==9'd262/*262:US*/) || (xpc10nz==9'd260/*260:US*/) || (xpc10nz==9'd258/*258:US*/) || 
              (xpc10nz==9'd256/*256:US*/) || (xpc10nz==8'd254/*254:US*/) || (xpc10nz==8'd252/*252:US*/) || (xpc10nz==8'd250/*250:US*/) || 
              (xpc10nz==8'd248/*248:US*/) || (xpc10nz==8'd246/*246:US*/) || (xpc10nz==8'd244/*244:US*/) || (xpc10nz==8'd242/*242:US*/) || 
              (xpc10nz==8'd240/*240:US*/) || (xpc10nz==8'd238/*238:US*/) || (xpc10nz==8'd236/*236:US*/) || (xpc10nz==8'd234/*234:US*/) || 
              (xpc10nz==8'd232/*232:US*/) || (xpc10nz==8'd230/*230:US*/) || (xpc10nz==8'd228/*228:US*/) || (xpc10nz==8'd226/*226:US*/) || 
              (xpc10nz==8'd224/*224:US*/) || (xpc10nz==8'd222/*222:US*/) || (xpc10nz==8'd220/*220:US*/) || (xpc10nz==8'd218/*218:US*/) || 
              (xpc10nz==8'd216/*216:US*/) || (xpc10nz==8'd214/*214:US*/) || (xpc10nz==8'd212/*212:US*/) || (xpc10nz==8'd210/*210:US*/) || 
              (xpc10nz==8'd208/*208:US*/) || (xpc10nz==8'd206/*206:US*/) || (xpc10nz==8'd204/*204:US*/) || (xpc10nz==8'd202/*202:US*/) || 
              (xpc10nz==8'd200/*200:US*/) || (xpc10nz==8'd198/*198:US*/) || (xpc10nz==8'd196/*196:US*/) || (xpc10nz==8'd194/*194:US*/) || 
              (xpc10nz==8'd192/*192:US*/) || (xpc10nz==8'd190/*190:US*/) || (xpc10nz==8'd188/*188:US*/) || (xpc10nz==8'd186/*186:US*/) || 
              (xpc10nz==8'd184/*184:US*/) || (xpc10nz==8'd182/*182:US*/) || (xpc10nz==8'd180/*180:US*/) || (xpc10nz==8'd178/*178:US*/) || 
              (xpc10nz==8'd176/*176:US*/) || (xpc10nz==8'd174/*174:US*/) || (xpc10nz==8'd172/*172:US*/) || (xpc10nz==8'd170/*170:US*/) || 
              (xpc10nz==8'd168/*168:US*/) || (xpc10nz==8'd166/*166:US*/) || (xpc10nz==8'd164/*164:US*/) || (xpc10nz==8'd162/*162:US*/) || 
              (xpc10nz==8'd160/*160:US*/) || (xpc10nz==8'd158/*158:US*/) || (xpc10nz==8'd156/*156:US*/) || (xpc10nz==8'd154/*154:US*/) || 
              (xpc10nz==8'd152/*152:US*/) || (xpc10nz==8'd150/*150:US*/) || (xpc10nz==8'd148/*148:US*/) || (xpc10nz==8'd146/*146:US*/) || 
              (xpc10nz==8'd144/*144:US*/) || (xpc10nz==8'd142/*142:US*/) || (xpc10nz==8'd140/*140:US*/) || (xpc10nz==8'd138/*138:US*/) || 
              (xpc10nz==8'd136/*136:US*/) || (xpc10nz==8'd134/*134:US*/) || (xpc10nz==8'd132/*132:US*/) || (xpc10nz==8'd130/*130:US*/) || 
              (xpc10nz==8'd128/*128:US*/) || (xpc10nz==7'd126/*126:US*/) || (xpc10nz==7'd124/*124:US*/) || (xpc10nz==7'd122/*122:US*/) || 
              (xpc10nz==7'd120/*120:US*/) || (xpc10nz==7'd118/*118:US*/) || (xpc10nz==7'd116/*116:US*/) || (xpc10nz==7'd114/*114:US*/) || 
              (xpc10nz==7'd112/*112:US*/) || (xpc10nz==7'd110/*110:US*/) || (xpc10nz==7'd108/*108:US*/) || (xpc10nz==7'd106/*106:US*/) || 
              (xpc10nz==7'd104/*104:US*/) || (xpc10nz==7'd102/*102:US*/) || (xpc10nz==7'd100/*100:US*/) || (xpc10nz==7'd98/*98:US*/) || 
              (xpc10nz==7'd96/*96:US*/) || (xpc10nz==7'd94/*94:US*/) || (xpc10nz==7'd92/*92:US*/) || (xpc10nz==7'd90/*90:US*/) || (xpc10nz
              ==7'd88/*88:US*/) || (xpc10nz==7'd86/*86:US*/) || (xpc10nz==7'd84/*84:US*/) || (xpc10nz==7'd82/*82:US*/) || (xpc10nz==7'd80
              /*80:US*/) || (xpc10nz==7'd78/*78:US*/) || (xpc10nz==7'd76/*76:US*/) || (xpc10nz==7'd74/*74:US*/) || (xpc10nz==7'd72/*72:US*/) || 
              (xpc10nz==7'd70/*70:US*/) || (xpc10nz==7'd68/*68:US*/) || (xpc10nz==7'd66/*66:US*/) || (xpc10nz==7'd64/*64:US*/) || (xpc10nz
              ==6'd62/*62:US*/) || (xpc10nz==6'd60/*60:US*/) || (xpc10nz==6'd58/*58:US*/) || (xpc10nz==6'd56/*56:US*/) || (xpc10nz==6'd54
              /*54:US*/) || (xpc10nz==6'd52/*52:US*/) || (xpc10nz==6'd50/*50:US*/) || (xpc10nz==6'd48/*48:US*/) || (xpc10nz==6'd46/*46:US*/) || 
              (xpc10nz==6'd44/*44:US*/) || (xpc10nz==6'd42/*42:US*/) || (xpc10nz==6'd40/*40:US*/) || (xpc10nz==6'd38/*38:US*/) || (xpc10nz
              ==6'd36/*36:US*/) || (xpc10nz==6'd34/*34:US*/) || (xpc10nz==6'd32/*32:US*/) || (xpc10nz==5'd30/*30:US*/) || (xpc10nz==5'd28
              /*28:US*/) || (xpc10nz==5'd26/*26:US*/) || (xpc10nz==5'd24/*24:US*/) || (xpc10nz==5'd22/*22:US*/) || (xpc10nz==5'd20/*20:US*/) || 
              (xpc10nz==5'd18/*18:US*/) || (xpc10nz==5'd16/*16:US*/) || (xpc10nz==4'd14/*14:US*/) || (xpc10nz==4'd12/*12:US*/) || (xpc10nz
              ==4'd10/*10:US*/) || (xpc10nz==4'd8/*8:US*/) || (xpc10nz==3'd6/*6:US*/) || (xpc10nz==3'd4/*4:US*/) || (xpc10nz==2'd2/*2:US*/) || 
              (xpc10nz==0/*0:US*/)? 1'd1: 1'd0);

               A_16_SS_CC_SCALbx10_ARA0_REN0 = ((xpc10nz==9'd409/*409:US*/)? 1'd1: 1'd0);
               A_64_SS_CC_SCALbx52_ARA0_WEN0 = ((xpc10nz==9'd407/*407:US*/) || (xpc10nz==9'd405/*405:US*/) || (xpc10nz==9'd414/*414:US*/)? 1'd1
              : 1'd0);

               A_SINT_CC_SCALbx16_ARA0_REN0 = ((xpc10nz==9'd418/*418:US*/)? 1'd1: 1'd0);
               A_64_SS_CC_SCALbx54_ARB0_WEN0 = (xpc10nz==9'd405/*405:US*/) || (xpc10nz==9'd407/*407:US*/) || (xpc10nz==9'd419/*419:US*/);
               A_64_SS_CC_SCALbx56_ARC0_REN0 = ((xpc10nz==9'd428/*428:US*/) || (xpc10nz==9'd432/*432:US*/)? 1'd1: 1'd0);
               A_64_SS_CC_SCALbx56_ARC0_WEN0 = (xpc10nz==9'd407/*407:US*/) || (xpc10nz==9'd405/*405:US*/) || ((64'hffffffffffffffff&64'h_ffff_ffff_ffff_fffe
              +A_64_SS_CC_SCALbx56_ARC0_RDD0)<A_64_SS_CC_SCALbx52_ARA0_RDD0) && (xpc10nz==9'd433/*433:US*/);

               A_64_SS_CC_SCALbx52_ARA0_REN0 = ((xpc10nz==9'd432/*432:US*/) || (xpc10nz==9'd438/*438:US*/)? 1'd1: 1'd0);
               A_64_SS_CC_SCALbx58_ARD0_REN0 = ((xpc10nz==9'd428/*428:US*/) || (xpc10nz==9'd438/*438:US*/)? 1'd1: 1'd0);
               A_64_SS_CC_SCALbx58_ARD0_WEN0 = (xpc10nz==9'd407/*407:US*/) || (xpc10nz==9'd405/*405:US*/) || ((64'hffffffffffffffff&64'h_ffff_ffff_ffff_fffe
              +A_64_SS_CC_SCALbx56_ARC0_RDD0)>=A_64_SS_CC_SCALbx52_ARA0_RDD0) && (xpc10nz==9'd433/*433:US*/) || (xpc10nz==9'd439/*439:US*/);

               A_64_SS_CC_SCALbx54_ARB0_REN0 = (xpc10nz==9'd424/*424:US*/) || (xpc10nz==9'd413/*413:US*/) || (xpc10nz==9'd444/*444:US*/) || 
              (TSPcr2_16_V_1<32'd77) && (xpc10nz==9'd461/*461:US*/);

               A_UINT_CC_SCALbx34_ARA0_REN0 = ((xpc10nz==9'd484/*484:US*/) || (xpc10nz==9'd482/*482:US*/) || (xpc10nz==9'd478/*478:US*/) || 
              (xpc10nz==9'd474/*474:US*/) || (xpc10nz==9'd457/*457:US*/) || (xpc10nz==9'd454/*454:US*/) || (xpc10nz==9'd451/*451:US*/) || 
              (xpc10nz==9'd448/*448:US*/) || (xpc10nz==9'd447/*447:US*/) || (xpc10nz==9'd450/*450:US*/) || (xpc10nz==9'd453/*453:US*/) || 
              (xpc10nz==9'd456/*456:US*/) || (xpc10nz==9'd473/*473:US*/) || (xpc10nz==9'd477/*477:US*/) || (xpc10nz==9'd481/*481:US*/) || 
              (xpc10nz==9'd487/*487:US*/)? 1'd1: 1'd0);

               A_SINT_CC_SCALbx26_ARJ0_WEN0 = (xpc10nz==9'd492/*492:US*/);
               A_16_SS_CC_SCALbx14_ARC0_REN0 = ((xpc10nz==9'd495/*495:US*/)? 1'd1: 1'd0);
               A_16_SS_CC_SCALbx12_ARB0_REN0 = ((xpc10nz==9'd409/*409:US*/) || (xpc10nz==9'd495/*495:US*/)? 1'd1: 1'd0);

              case (xpc10nz)
                  0/*0:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_b2f7_40b4;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd255;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd10;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd399;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd108;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd74;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd110;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd76;
                       A_16_SS_CC_SCALbx12_ARB0_WRD0 = 16'd121;
                       A_16_SS_CC_SCALbx12_ARB0_AD0 = 6'd19;
                       end 
                      
                  1'd1/*1:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_b636_5d03;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd254;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd398;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd112;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd73;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd101;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd75;
                       A_16_SS_CC_SCALbx12_ARB0_WRD0 = 16'd119;
                       A_16_SS_CC_SCALbx12_ARB0_AD0 = 6'd18;
                       end 
                      
                  2'd2/*2:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_b975_7bda;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd253;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd397;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd105;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd72;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd113;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd74;
                       A_16_SS_CC_SCALbx12_ARB0_WRD0 = 16'd118;
                       A_16_SS_CC_SCALbx12_ARB0_AD0 = 6'd17;
                       end 
                      
                  2'd3/*3:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_bdb4_666d;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd252;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffd;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd396;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd116;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd71;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd114;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd73;
                       A_16_SS_CC_SCALbx12_ARB0_WRD0 = 16'd116;
                       A_16_SS_CC_SCALbx12_ARB0_AD0 = 6'd16;
                       end 
                      
                  3'd4/*4:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_a3f3_3668;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd251;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffd;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd395;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd101;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd70;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd118;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd72;
                       A_16_SS_CC_SCALbx12_ARB0_WRD0 = 16'd115;
                       A_16_SS_CC_SCALbx12_ARB0_AD0 = 6'd15;
                       end 
                      
                  3'd5/*5:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_a732_2bdf;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd250;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffc;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd394;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd121;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd69;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd101;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd71;
                       A_16_SS_CC_SCALbx12_ARB0_WRD0 = 16'd114;
                       A_16_SS_CC_SCALbx12_ARB0_AD0 = 6'd14;
                       end 
                      
                  3'd6/*6:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_ac71_0d06;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd249;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffc;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd393;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd103;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd68;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd107;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd70;
                       A_16_SS_CC_SCALbx12_ARB0_WRD0 = 16'd113;
                       A_16_SS_CC_SCALbx12_ARB0_AD0 = 6'd13;
                       end 
                      
                  3'd7/*7:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_b0b0_10b1;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd248;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffb;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd392;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd113;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd67;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd97;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd69;
                       A_16_SS_CC_SCALbx12_ARB0_WRD0 = 16'd112;
                       A_16_SS_CC_SCALbx12_ARB0_AD0 = 6'd12;
                       end 
                      
                  4'd8/*8:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_98ff_ad0c;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd247;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd391;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd105;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd66;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd101;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd68;
                       A_16_SS_CC_SCALbx12_ARB0_WRD0 = 16'd110;
                       A_16_SS_CC_SCALbx12_ARB0_AD0 = 6'd11;
                       end 
                      
                  4'd9/*9:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_943e_b0bb;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd246;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd390;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd114;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd65;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd101;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd67;
                       A_16_SS_CC_SCALbx12_ARB0_WRD0 = 16'd109;
                       A_16_SS_CC_SCALbx12_ARB0_AD0 = 6'd10;
                       end 
                      
                  4'd10/*10:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_9f7d_9662;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd245;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_ffff;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd389;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd97;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd64;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd108;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd66;
                       A_16_SS_CC_SCALbx12_ARB0_WRD0 = 16'd108;
                       A_16_SS_CC_SCALbx12_ARB0_AD0 = 6'd9;
                       end 
                      
                  4'd11/*11:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_9bbc_8bd5;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd244;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffc;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd388;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd118;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd63;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd97;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd65;
                       A_16_SS_CC_SCALbx12_ARB0_WRD0 = 16'd107;
                       A_16_SS_CC_SCALbx12_ARB0_AD0 = 6'd8;
                       end 
                      
                  4'd12/*12:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_85fb_dbd0;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd243;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_ffff;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd387;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd101;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd62;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd101;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd64;
                       A_16_SS_CC_SCALbx12_ARB0_WRD0 = 16'd105;
                       A_16_SS_CC_SCALbx12_ARB0_AD0 = 6'd7;
                       end 
                      
                  4'd13/*13:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_813a_c667;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd242;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd386;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd101;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd61;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd113;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd63;
                       A_16_SS_CC_SCALbx12_ARB0_WRD0 = 16'd104;
                       A_16_SS_CC_SCALbx12_ARB0_AD0 = 6'd6;
                       end 
                      
                  4'd14/*14:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_8e79_e0be;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd241;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffb;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd385;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd118;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd60;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd115;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd62;
                       A_16_SS_CC_SCALbx12_ARB0_WRD0 = 16'd103;
                       A_16_SS_CC_SCALbx12_ARB0_AD0 = 6'd5;
                       end 
                      
                  4'd15/*15:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_8ab8_fd09;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd240;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd7;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd384;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd108;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd59;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd103;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd61;
                       A_16_SS_CC_SCALbx12_ARB0_WRD0 = 16'd102;
                       A_16_SS_CC_SCALbx12_ARB0_AD0 = 6'd4;
                       end 
                      
                  5'd16/*16:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_fee6_9bc4;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd239;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffc;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd383;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd100;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd58;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd119;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd60;
                       A_16_SS_CC_SCALbx12_ARB0_WRD0 = 16'd101;
                       A_16_SS_CC_SCALbx12_ARB0_AD0 = 6'd3;
                       end 
                      
                  5'd17/*17:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_fa27_8673;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd238;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffc;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd382;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd101;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd57;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd118;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd59;
                       A_16_SS_CC_SCALbx12_ARB0_WRD0 = 16'd100;
                       A_16_SS_CC_SCALbx12_ARB0_AD0 = 6'd2;
                       end 
                      
                  5'd18/*18:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_f564_a0aa;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd237;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd381;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd101;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd56;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd101;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd58;
                       A_16_SS_CC_SCALbx12_ARB0_WRD0 = 16'd99;
                       A_16_SS_CC_SCALbx12_ARB0_AD0 = 6'd1;
                       end 
                      
                  5'd19/*19:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_f1a5_bd1d;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd236;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffd;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd380;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd108;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd55;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd108;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd57;
                       A_16_SS_CC_SCALbx12_ARB0_WRD0 = 16'd97;
                       A_16_SS_CC_SCALbx12_ARB0_AD0 = 6'd0;
                       end 
                      
                  5'd20/*20:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_efe2_ed18;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd235;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd379;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd114;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd54;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd115;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd56;
                       end 
                      
                  5'd21/*21:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_eb23_f0af;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd234;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd17;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd378;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd108;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd53;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd114;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd55;
                       end 
                      
                  5'd22/*22:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_e860_d676;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd233;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffa;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd377;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd100;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd52;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd107;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd54;
                       end 
                      
                  5'd23/*23:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_e4a1_cbc1;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd232;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffb;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd376;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd108;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd51;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd118;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd53;
                       end 
                      
                  5'd24/*24:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_dcee_767c;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd231;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd375;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd114;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd50;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd105;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd52;
                       end 
                      
                  5'd25/*25:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_e02f_6bcb;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd230;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd2;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd374;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd104;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd49;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd113;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd51;
                       end 
                      
                  5'd26/*26:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_d36c_4d12;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd229;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffb;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd373;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd115;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd48;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd108;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd50;
                       end 
                      
                  5'd27/*27:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_d7ad_50a5;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd228;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffa;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd372;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd112;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd47;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd107;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd49;
                       end 
                      
                  5'd28/*28:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_c9ea_00a0;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd227;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffc;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd371;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd112;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd46;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd108;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd48;
                       end 
                      
                  5'd29/*29:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_cd2b_1d17;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd226;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffc;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd370;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd116;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd45;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd121;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd47;
                       end 
                      
                  5'd30/*30:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_c268_3bce;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd225;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd369;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd118;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd44;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd108;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd46;
                       end 
                      
                  5'd31/*31:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_c6a9_2679;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd224;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffd;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd368;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd114;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd43;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd107;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd45;
                       end 
                      
                  6'd32/*32:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_29d4_f654;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd223;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffb;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd367;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd121;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd42;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd109;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd44;
                       end 
                      
                  6'd33/*33:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_2d15_ebe3;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd222;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffd;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd366;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd116;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd41;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd100;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd43;
                       end 
                      
                  6'd34/*34:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_2056_cd3a;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd221;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fff9;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd365;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd112;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd40;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd103;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd42;
                       end 
                      
                  6'd35/*35:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_2497_d08d;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd220;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd364;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd103;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd39;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd119;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd41;
                       end 
                      
                  6'd36/*36:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_3ad0_8088;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd219;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fff9;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd363;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd101;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd38;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd113;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd40;
                       end 
                      
                  6'd37/*37:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_3e11_9d3f;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd218;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fff9;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd362;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd103;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd37;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd115;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd39;
                       end 
                      
                  6'd38/*38:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_3352_bbe6;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd217;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fff8;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd361;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd101;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd36;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd104;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd38;
                       end 
                      
                  6'd39/*39:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_3793_a651;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd216;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffa;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd360;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd118;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd35;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd104;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd37;
                       end 
                      
                  6'd40/*40:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'hfdc_1bec;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd215;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd359;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd114;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd34;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd112;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd36;
                       end 
                      
                  6'd41/*41:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'hb1d_065b;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd214;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffa;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd358;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd99;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd33;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd110;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd35;
                       end 
                      
                  6'd42/*42:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h65e_2082;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd213;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd4;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd357;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd103;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd32;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd107;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd34;
                       end 
                      
                  6'd43/*43:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h29f_3d35;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd212;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd356;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd108;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd31;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd107;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd33;
                       end 
                      
                  6'd44/*44:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_1cd8_6d30;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd211;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_ffff;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd355;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd114;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd30;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd118;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd32;
                       end 
                      
                  6'd45/*45:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_1819_7087;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd210;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd354;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd107;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd29;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd105;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd31;
                       end 
                      
                  6'd46/*46:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_155a_565e;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd209;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd353;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd108;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd28;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd102;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd30;
                       end 
                      
                  6'd47/*47:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_119b_4be9;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd208;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_ffff;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd352;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd105;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd27;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd107;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd29;
                       end 
                      
                  6'd48/*48:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_65c5_2d24;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd207;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd351;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd97;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd26;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd108;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd28;
                       end 
                      
                  6'd49/*49:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_6104_3093;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd206;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd2;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd350;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd105;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd25;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd112;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd27;
                       end 
                      
                  6'd50/*50:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_6c47_164a;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd205;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd2;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd349;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd113;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd24;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd112;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd26;
                       end 
                      
                  6'd51/*51:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_6886_0bfd;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd204;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd348;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd101;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd23;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd101;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd25;
                       end 
                      
                  6'd52/*52:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_76c1_5bf8;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd203;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd4;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd347;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd97;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd22;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd114;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd24;
                       end 
                      
                  6'd53/*53:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_7200_464f;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd202;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd346;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd101;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd21;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd107;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd23;
                       end 
                      
                  6'd54/*54:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_7f43_6096;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd201;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_ffff;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd345;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd112;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd20;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd101;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd22;
                       end 
                      
                  6'd55/*55:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_7b82_7d21;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd200;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_ffff;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd344;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd121;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd19;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd108;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd21;
                       end 
                      
                  6'd56/*56:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_43cd_c09c;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd199;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd343;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd115;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd18;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd100;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd20;
                       end 
                      
                  6'd57/*57:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_470c_dd2b;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd198;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd342;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd116;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd17;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd99;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd19;
                       end 
                      
                  6'd58/*58:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_4a4f_fbf2;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd197;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd341;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd103;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd16;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd100;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd18;
                       end 
                      
                  6'd59/*59:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_4e8e_e645;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd196;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd340;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd108;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd15;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd107;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd17;
                       end 
                      
                  6'd60/*60:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_50c9_b640;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd195;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffd;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd339;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd108;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd14;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd108;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd16;
                       end 
                      
                  6'd61/*61:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_5408_abf7;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd194;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffb;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd338;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd114;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd13;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd108;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd15;
                       end 
                      
                  6'd62/*62:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_594b_8d2e;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd193;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd337;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd110;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd12;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd121;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd14;
                       end 
                      
                  6'd63/*63:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_5d8a_9099;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd192;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd3;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd336;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd97;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd11;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd101;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd13;
                       end 
                      
                  7'd64/*64:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_8671_30c3;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd191;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd1;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd335;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd121;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd10;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd113;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd12;
                       end 
                      
                  7'd65/*65:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_82b0_2d74;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd190;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_ffff;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd334;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd101;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd9;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd107;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd11;
                       end 
                      
                  7'd66/*66:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_8df3_0bad;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd189;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_ffff;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd333;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd112;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd8;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd97;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd10;
                       end 
                      
                  7'd67/*67:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_8932_161a;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd188;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd332;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd114;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd7;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd101;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd9;
                       end 
                      
                  7'd68/*68:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_9775_461f;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd187;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd331;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd102;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd6;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd116;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd8;
                       end 
                      
                  7'd69/*69:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_93b4_5ba8;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd186;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_ffff;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd330;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd112;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd5;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd107;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd7;
                       end 
                      
                  7'd70/*70:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_a0f7_7d71;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd185;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd329;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd105;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd4;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd116;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd6;
                       end 
                      
                  7'd71/*71:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_9c36_60c6;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd184;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd328;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd97;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd3;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd105;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd5;
                       end 
                      
                  7'd72/*72:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_a479_dd7b;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd183;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd327;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd101;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd2;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd108;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd4;
                       end 
                      
                  7'd73/*73:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_a8b8_c0cc;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd182;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_ffff;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd326;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd112;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd1;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd107;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd3;
                       end 
                      
                  7'd74/*74:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_abfb_e615;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd181;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd325;
                       A_16_SS_CC_SCALbx10_ARA0_WRD0 = 16'd112;
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = 8'd0;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd104;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd2;
                       end 
                      
                  7'd75/*75:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_af3a_fba2;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd180;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffd;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd324;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd107;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd1;
                       end 
                      
                  7'd76/*76:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_b17d_aba7;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd179;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd323;
                       A_16_SS_CC_SCALbx14_ARC0_WRD0 = 16'd100;
                       A_16_SS_CC_SCALbx14_ARC0_AD0 = 8'd0;
                       end 
                      
                  7'd77/*77:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_b5bc_b610;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd178;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd322;
                       end 
                      
                  7'd78/*78:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_baff_90c9;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd177;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd321;
                       end 
                      
                  7'd79/*79:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_be3e_8d7e;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd176;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd1;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd320;
                       end 
                      
                  7'd80/*80:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_ca60_ebb3;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd175;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffd;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd319;
                       end 
                      
                  7'd81/*81:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_cea1_f604;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd174;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd318;
                       end 
                      
                  7'd82/*82:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_c1e2_d0dd;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd173;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_ffff;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd317;
                       end 
                      
                  7'd83/*83:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_c523_cd6a;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd172;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd1;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd316;
                       end 
                      
                  7'd84/*84:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_db64_9d6f;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd171;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd2;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd315;
                       end 
                      
                  7'd85/*85:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_dfa5_80d8;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd170;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd314;
                       end 
                      
                  7'd86/*86:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_d4e6_a601;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd169;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_ffff;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd313;
                       end 
                      
                  7'd87/*87:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_d827_bbb6;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd168;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd1;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd312;
                       end 
                      
                  7'd88/*88:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_f068_060b;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd167;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd1;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd311;
                       end 
                      
                  7'd89/*89:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_eca9_1bbc;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd166;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd310;
                       end 
                      
                  7'd90/*90:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_e7ea_3d65;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd165;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffd;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd309;
                       end 
                      
                  7'd91/*91:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_e32b_20d2;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd164;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd308;
                       end 
                      
                  7'd92/*92:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_fd6c_70d7;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd163;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_ffff;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd307;
                       end 
                      
                  7'd93/*93:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_f9ad_6d60;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd162;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_ffff;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd306;
                       end 
                      
                  7'd94/*94:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_f6ee_4bb9;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd161;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd1;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd305;
                       end 
                      
                  7'd95/*95:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_f22f_560e;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd160;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffd;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd304;
                       end 
                      
                  7'd96/*96:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_1d52_8623;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd159;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd303;
                       end 
                      
                  7'd97/*97:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_1993_9b94;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd158;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd302;
                       end 
                      
                  7'd98/*98:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_14d0_bd4d;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd157;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd301;
                       end 
                      
                  7'd99/*99:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_1011_a0fa;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd156;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd1;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd300;
                       end 
                      
                  7'd100/*100:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'he56_f0ff;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd155;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffc;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd299;
                       end 
                      
                  7'd101/*101:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'ha97_ed48;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd154;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd2;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd298;
                       end 
                      
                  7'd102/*102:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h7d4_cb91;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd153;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd297;
                       end 
                      
                  7'd103/*103:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h315_d626;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd152;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_ffff;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd296;
                       end 
                      
                  7'd104/*104:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_3b5a_6b9b;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd151;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd295;
                       end 
                      
                  7'd105/*105:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_3f9b_762c;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd150;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd6;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd294;
                       end 
                      
                  7'd106/*106:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_32d8_50f5;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd149;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd1;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd293;
                       end 
                      
                  7'd107/*107:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_3619_4d42;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd148;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd292;
                       end 
                      
                  7'd108/*108:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_285e_1d47;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd147;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd291;
                       end 
                      
                  7'd109/*109:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_2c9f_00f0;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd146;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd290;
                       end 
                      
                  7'd110/*110:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_21dc_2629;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd145;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffd;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd289;
                       end 
                      
                  7'd111/*111:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_251d_3b9e;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd144;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd3;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd288;
                       end 
                      
                  7'd112/*112:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_5143_5d53;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd143;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd287;
                       end 
                      
                  7'd113/*113:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_5582_40e4;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd142;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd2;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd286;
                       end 
                      
                  7'd114/*114:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_58c1_663d;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd141;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffd;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd285;
                       end 
                      
                  7'd115/*115:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_5c00_7b8a;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd140;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffc;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd284;
                       end 
                      
                  7'd116/*116:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_4247_2b8f;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd139;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_ffff;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd283;
                       end 
                      
                  7'd117/*117:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_4686_3638;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd138;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_ffff;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd282;
                       end 
                      
                  7'd118/*118:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_4bc5_10e1;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd137;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffc;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd281;
                       end 
                      
                  7'd119/*119:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_4f04_0d56;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd136;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd280;
                       end 
                      
                  7'd120/*120:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_774b_b0eb;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd135;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffc;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd279;
                       end 
                      
                  7'd121/*121:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_738a_ad5c;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd134;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffb;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd278;
                       end 
                      
                  7'd122/*122:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_7ec9_8b85;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd133;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd277;
                       end 
                      
                  7'd123/*123:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_7a08_9632;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd132;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_ffff;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd276;
                       end 
                      
                  7'd124/*124:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_644f_c637;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd131;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_ffff;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd275;
                       end 
                      
                  7'd125/*125:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_608e_db80;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd130;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd1;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd274;
                       end 
                      
                  7'd126/*126:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_6dcd_fd59;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd129;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd4;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd273;
                       end 
                      
                  7'd127/*127:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_690c_e0ee;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd128;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd272;
                       end 
                      
                  8'd128/*128:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_d9fb_a05a;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd127;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd1;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd271;
                       end 
                      
                  8'd129/*129:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_dd3a_bded;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd126;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_ffff;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd270;
                       end 
                      
                  8'd130/*130:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_d279_9b34;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd125;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd269;
                       end 
                      
                  8'd131/*131:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_d6b8_8683;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd124;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd1;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd268;
                       end 
                      
                  8'd132/*132:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_ccff_d686;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd123;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd267;
                       end 
                      
                  8'd133/*133:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_d03e_cb31;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd122;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd3;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd266;
                       end 
                      
                  8'd134/*134:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_c37d_ede8;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd121;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_ffff;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd265;
                       end 
                      
                  8'd135/*135:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_c7bc_f05f;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd120;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffb;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd264;
                       end 
                      
                  8'd136/*136:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_fff3_4de2;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd119;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd2;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd263;
                       end 
                      
                  8'd137/*137:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_fb32_5055;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd118;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd2;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd262;
                       end 
                      
                  8'd138/*138:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_f871_768c;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd117;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffb;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd261;
                       end 
                      
                  8'd139/*139:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_f4b0_6b3b;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd116;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd260;
                       end 
                      
                  8'd140/*140:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_eef7_3b3e;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd115;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffb;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd259;
                       end 
                      
                  8'd141/*141:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_ea36_2689;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd114;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffa;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd258;
                       end 
                      
                  8'd142/*142:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_e575_0050;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd113;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_ffff;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd257;
                       end 
                      
                  8'd143/*143:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_e1b4_1de7;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd112;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd256;
                       end 
                      
                  8'd144/*144:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_95ea_7b2a;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd111;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd1;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd255;
                       end 
                      
                  8'd145/*145:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_912b_669d;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd110;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd254;
                       end 
                      
                  8'd146/*146:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_9e68_4044;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd109;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd253;
                       end 
                      
                  8'd147/*147:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_9aa9_5df3;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd108;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd6;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd252;
                       end 
                      
                  8'd148/*148:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_88ee_0df6;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd107;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_ffff;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd251;
                       end 
                      
                  8'd149/*149:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_842f_1041;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd106;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd250;
                       end 
                      
                  8'd150/*150:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_8f6c_3698;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd105;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffd;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd249;
                       end 
                      
                  8'd151/*151:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_8bad_2b2f;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd104;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_ffff;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd248;
                       end 
                      
                  8'd152/*152:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_b3e2_9692;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd103;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd247;
                       end 
                      
                  8'd153/*153:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_b723_8b25;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd102;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd246;
                       end 
                      
                  8'd154/*154:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_bc60_adfc;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd101;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_ffff;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd245;
                       end 
                      
                  8'd155/*155:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_c0a1_b04b;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd100;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffb;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd244;
                       end 
                      
                  8'd156/*156:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_a2e6_e04e;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd99;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_ffff;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd243;
                       end 
                      
                  8'd157/*157:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_a627_fdf9;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd98;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_ffff;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd242;
                       end 
                      
                  8'd158/*158:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_a964_db20;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd97;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffd;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd241;
                       end 
                      
                  8'd159/*159:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_ada5_c697;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd96;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd1;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd240;
                       end 
                      
                  8'd160/*160:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_40d8_16ba;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd95;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd239;
                       end 
                      
                  8'd161/*161:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_4419_0b0d;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd94;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffc;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd238;
                       end 
                      
                  8'd162/*162:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_495a_2dd4;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd93;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd237;
                       end 
                      
                  8'd163/*163:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_4d9b_3063;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd92;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd236;
                       end 
                      
                  8'd164/*164:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_53dc_6066;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd91;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd1;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd235;
                       end 
                      
                  8'd165/*165:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_571d_7dd1;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd90;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd234;
                       end 
                      
                  8'd166/*166:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_5a5e_5b08;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd89;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd1;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd233;
                       end 
                      
                  8'd167/*167:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_5e9f_46bf;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd88;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_ffff;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd232;
                       end 
                      
                  8'd168/*168:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_66d0_fb02;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd87;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd2;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd231;
                       end 
                      
                  8'd169/*169:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_6211_e6b5;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd86;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd230;
                       end 
                      
                  8'd170/*170:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_6f52_c06c;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd85;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffd;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd229;
                       end 
                      
                  8'd171/*171:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_6b93_dddb;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd84;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd1;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd228;
                       end 
                      
                  8'd172/*172:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_75d4_8dde;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd83;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd227;
                       end 
                      
                  8'd173/*173:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_7115_9069;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd82;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd2;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd226;
                       end 
                      
                  8'd174/*174:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_7c56_b6b0;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd81;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd225;
                       end 
                      
                  8'd175/*175:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_7897_ab07;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd80;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffc;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd224;
                       end 
                      
                  8'd176/*176:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'hcc9_cdca;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd79;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd1;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd223;
                       end 
                      
                  8'd177/*177:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h808_d07d;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd78;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd2;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd222;
                       end 
                      
                  8'd178/*178:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h54b_f6a4;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd77;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffc;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd221;
                       end 
                      
                  8'd179/*179:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h18a_eb13;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd76;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd220;
                       end 
                      
                  8'd180/*180:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_1fcd_bb16;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd75;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd219;
                       end 
                      
                  8'd181/*181:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_1b0c_a6a1;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd74;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffc;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd218;
                       end 
                      
                  8'd182/*182:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_164f_8078;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd73;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd2;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd217;
                       end 
                      
                  8'd183/*183:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_128e_9dcf;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd72;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_ffff;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd216;
                       end 
                      
                  8'd184/*184:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_2ac1_2072;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd71;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd215;
                       end 
                      
                  8'd185/*185:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_2e00_3dc5;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd70;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd214;
                       end 
                      
                  8'd186/*186:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_2343_1b1c;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd69;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_ffff;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd213;
                       end 
                      
                  8'd187/*187:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_2782_06ab;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd68;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd212;
                       end 
                      
                  8'd188/*188:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_39c5_56ae;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd67;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd211;
                       end 
                      
                  8'd189/*189:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_3d04_4b19;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd66;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd6;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd210;
                       end 
                      
                  8'd190/*190:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_3047_6dc0;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd65;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd4;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd209;
                       end 
                      
                  8'd191/*191:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_3486_7077;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd64;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd208;
                       end 
                      
                  8'd192/*192:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_ed7d_d02d;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd63;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd2;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd207;
                       end 
                      
                  8'd193/*193:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_e9bc_cd9a;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd62;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd206;
                       end 
                      
                  8'd194/*194:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_e6ff_eb43;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd61;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffd;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd205;
                       end 
                      
                  8'd195/*195:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_e23e_f6f4;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd60;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd204;
                       end 
                      
                  8'd196/*196:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_ff79_a6f1;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd59;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd203;
                       end 
                      
                  8'd197/*197:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_fcb8_bb46;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd58;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffd;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd202;
                       end 
                      
                  8'd198/*198:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_f7fb_9d9f;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd57;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffb;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd201;
                       end 
                      
                  8'd199/*199:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_f33a_8028;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd56;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_ffff;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd200;
                       end 
                      
                  8'd200/*200:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_cb75_3d95;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd55;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_ffff;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd199;
                       end 
                      
                  8'd201/*201:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_cfb4_2022;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd54;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd198;
                       end 
                      
                  8'd202/*202:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_c4f7_06fb;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd53;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd2;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd197;
                       end 
                      
                  8'd203/*203:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_c836_1b4c;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd52;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd196;
                       end 
                      
                  8'd204/*204:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_da71_4b49;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd51;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffd;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd195;
                       end 
                      
                  8'd205/*205:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_deb0_56fe;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd50;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffd;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd194;
                       end 
                      
                  8'd206/*206:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_d1f3_7027;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd49;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd193;
                       end 
                      
                  8'd207/*207:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_d532_6d90;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd48;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffd;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd192;
                       end 
                      
                  8'd208/*208:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_a16c_0b5d;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd47;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffd;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd191;
                       end 
                      
                  8'd209/*209:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_a5ad_16ea;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd46;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd4;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd190;
                       end 
                      
                  8'd210/*210:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_aaee_3033;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd45;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd6;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd189;
                       end 
                      
                  8'd211/*211:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_ae2f_2d84;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd44;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffd;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd188;
                       end 
                      
                  8'd212/*212:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_b468_7d81;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd43;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd2;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd187;
                       end 
                      
                  8'd213/*213:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_b8a9_6036;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd42;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd186;
                       end 
                      
                  8'd214/*214:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_bbea_46ef;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd41;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffc;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd185;
                       end 
                      
                  8'd215/*215:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_bf2b_5b58;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd40;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd2;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd184;
                       end 
                      
                  8'd216/*216:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_8764_e6e5;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd39;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffd;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd183;
                       end 
                      
                  8'd217/*217:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_83a5_fb52;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd38;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffc;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd182;
                       end 
                      
                  8'd218/*218:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_90e6_dd8b;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd37;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffa;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd181;
                       end 
                      
                  8'd219/*219:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_8c27_c03c;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd36;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd180;
                       end 
                      
                  8'd220/*220:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_9660_9039;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd35;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffc;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd179;
                       end 
                      
                  8'd221/*221:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_92a1_8d8e;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd34;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffd;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd178;
                       end 
                      
                  8'd222/*222:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_9de2_ab57;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd33;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd177;
                       end 
                      
                  8'd223/*223:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_9923_b6e0;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd32;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd176;
                       end 
                      
                  8'd224/*224:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_745e_66cd;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd31;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd175;
                       end 
                      
                  8'd225/*225:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_709f_7b7a;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd30;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd3;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd174;
                       end 
                      
                  8'd226/*226:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_7ddc_5da3;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd29;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd1;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd173;
                       end 
                      
                  8'd227/*227:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_791d_4014;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd28;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_ffff;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd172;
                       end 
                      
                  8'd228/*228:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_675a_1011;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd27;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd1;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd171;
                       end 
                      
                  8'd229/*229:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_639b_0da6;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd26;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd170;
                       end 
                      
                  8'd230/*230:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_6ed8_2b7f;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd25;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffd;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd169;
                       end 
                      
                  8'd231/*231:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_6a19_36c8;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd24;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd5;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd168;
                       end 
                      
                  8'd232/*232:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_5256_8b75;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd23;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd167;
                       end 
                      
                  8'd233/*233:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_5697_96c2;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd22;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd166;
                       end 
                      
                  8'd234/*234:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_5bd4_b01b;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd21;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd165;
                       end 
                      
                  8'd235/*235:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_5f15_adac;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd20;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffb;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd164;
                       end 
                      
                  8'd236/*236:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_4152_fda9;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd19;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd163;
                       end 
                      
                  8'd237/*237:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_4593_e01e;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd18;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd162;
                       end 
                      
                  8'd238/*238:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_48d0_c6c7;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd17;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffb;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd161;
                       end 
                      
                  8'd239/*239:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_4c11_db70;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd16;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_ffff;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd160;
                       end 
                      
                  8'd240/*240:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_384f_bdbd;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd15;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_ffff;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd159;
                       end 
                      
                  8'd241/*241:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_3c8e_a00a;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd14;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffb;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd158;
                       end 
                      
                  8'd242/*242:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_31cd_86d3;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd13;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd4;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd157;
                       end 
                      
                  8'd243/*243:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_350c_9b64;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd12;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd156;
                       end 
                      
                  8'd244/*244:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_2b4b_cb61;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd11;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_ffff;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd155;
                       end 
                      
                  8'd245/*245:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_2f8a_d6d6;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd10;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd154;
                       end 
                      
                  8'd246/*246:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_22c9_f00f;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd9;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd153;
                       end 
                      
                  8'd247/*247:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_2608_edb8;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd8;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd152;
                       end 
                      
                  8'd248/*248:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_1e47_5005;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd7;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd151;
                       end 
                      
                  8'd249/*249:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_1a86_4db2;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd6;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd2;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd150;
                       end 
                      
                  8'd250/*250:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_17c5_6b6b;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd5;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd2;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd149;
                       end 
                      
                  8'd251/*251:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h_1304_76dc;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd4;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd148;
                       end 
                      
                  8'd252/*252:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'hd43_26d9;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd3;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd5;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd147;
                       end 
                      
                  8'd253/*253:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h982_3b6e;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd2;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd146;
                       end 
                      
                  8'd254/*254:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'h4c1_1db7;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd1;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffd;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd145;
                       end 
                      
                  8'd255/*255:US*/:  begin 
                       A_UINT_CC_SCALbx34_ARA0_WRD0 = 32'd0;
                       A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd0;
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd1;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd144;
                       end 
                      
                  9'd256/*256:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd143;
                       end 
                      
                  9'd257/*257:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd142;
                       end 
                      
                  9'd258/*258:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd141;
                       end 
                      
                  9'd259/*259:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_ffff;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd140;
                       end 
                      
                  9'd260/*260:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd139;
                       end 
                      
                  9'd261/*261:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffd;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd138;
                       end 
                      
                  9'd262/*262:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd137;
                       end 
                      
                  9'd263/*263:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_ffff;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd136;
                       end 
                      
                  9'd264/*264:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_ffff;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd135;
                       end 
                      
                  9'd265/*265:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd2;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd134;
                       end 
                      
                  9'd266/*266:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd3;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd133;
                       end 
                      
                  9'd267/*267:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd132;
                       end 
                      
                  9'd268/*268:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd2;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd131;
                       end 
                      
                  9'd269/*269:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd130;
                       end 
                      
                  9'd270/*270:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd129;
                       end 
                      
                  9'd271/*271:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd128;
                       end 
                      
                  9'd272/*272:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd127;
                       end 
                      
                  9'd273/*273:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd6;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd126;
                       end 
                      
                  9'd274/*274:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd125;
                       end 
                      
                  9'd275/*275:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd124;
                       end 
                      
                  9'd276/*276:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd1;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd123;
                       end 
                      
                  9'd277/*277:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd1;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd122;
                       end 
                      
                  9'd278/*278:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffd;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd121;
                       end 
                      
                  9'd279/*279:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_ffff;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd120;
                       end 
                      
                  9'd280/*280:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffb;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd119;
                       end 
                      
                  9'd281/*281:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fff9;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd118;
                       end 
                      
                  9'd282/*282:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_ffff;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd117;
                       end 
                      
                  9'd283/*283:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd116;
                       end 
                      
                  9'd284/*284:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd1;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd115;
                       end 
                      
                  9'd285/*285:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffd;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd114;
                       end 
                      
                  9'd286/*286:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_ffff;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd113;
                       end 
                      
                  9'd287/*287:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_ffff;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd112;
                       end 
                      
                  9'd288/*288:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd111;
                       end 
                      
                  9'd289/*289:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffd;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd110;
                       end 
                      
                  9'd290/*290:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffc;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd109;
                       end 
                      
                  9'd291/*291:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd108;
                       end 
                      
                  9'd292/*292:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffd;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd107;
                       end 
                      
                  9'd293/*293:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd106;
                       end 
                      
                  9'd294/*294:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd5;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd105;
                       end 
                      
                  9'd295/*295:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffb;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd104;
                       end 
                      
                  9'd296/*296:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd103;
                       end 
                      
                  9'd297/*297:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd1;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd102;
                       end 
                      
                  9'd298/*298:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffd;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd101;
                       end 
                      
                  9'd299/*299:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd1;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd100;
                       end 
                      
                  9'd300/*300:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd7;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd99;
                       end 
                      
                  9'd301/*301:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd98;
                       end 
                      
                  9'd302/*302:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_ffff;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd97;
                       end 
                      
                  9'd303/*303:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffd;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd96;
                       end 
                      
                  9'd304/*304:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffd;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd95;
                       end 
                      
                  9'd305/*305:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffc;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd94;
                       end 
                      
                  9'd306/*306:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffb;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd93;
                       end 
                      
                  9'd307/*307:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffb;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd92;
                       end 
                      
                  9'd308/*308:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffc;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd91;
                       end 
                      
                  9'd309/*309:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd90;
                       end 
                      
                  9'd310/*310:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd2;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd89;
                       end 
                      
                  9'd311/*311:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffb;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd88;
                       end 
                      
                  9'd312/*312:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd1;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd87;
                       end 
                      
                  9'd313/*313:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd86;
                       end 
                      
                  9'd314/*314:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffb;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd85;
                       end 
                      
                  9'd315/*315:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd9;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd84;
                       end 
                      
                  9'd316/*316:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffb;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd83;
                       end 
                      
                  9'd317/*317:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffa;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd82;
                       end 
                      
                  9'd318/*318:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffc;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd81;
                       end 
                      
                  9'd319/*319:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffc;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd80;
                       end 
                      
                  9'd320/*320:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffc;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd79;
                       end 
                      
                  9'd321/*321:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fff9;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd78;
                       end 
                      
                  9'd322/*322:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd77;
                       end 
                      
                  9'd323/*323:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd76;
                       end 
                      
                  9'd324/*324:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd75;
                       end 
                      
                  9'd325/*325:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_ffff;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd74;
                       end 
                      
                  9'd326/*326:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd2;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd73;
                       end 
                      
                  9'd327/*327:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_ffff;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd72;
                       end 
                      
                  9'd328/*328:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd1;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd71;
                       end 
                      
                  9'd329/*329:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd70;
                       end 
                      
                  9'd330/*330:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffd;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd69;
                       end 
                      
                  9'd331/*331:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd68;
                       end 
                      
                  9'd332/*332:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd67;
                       end 
                      
                  9'd333/*333:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd1;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd66;
                       end 
                      
                  9'd334/*334:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd65;
                       end 
                      
                  9'd335/*335:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffb;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd64;
                       end 
                      
                  9'd336/*336:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd4;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd63;
                       end 
                      
                  9'd337/*337:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd3;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd62;
                       end 
                      
                  9'd338/*338:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffb;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd61;
                       end 
                      
                  9'd339/*339:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd60;
                       end 
                      
                  9'd340/*340:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffc;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd59;
                       end 
                      
                  9'd341/*341:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fff9;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd58;
                       end 
                      
                  9'd342/*342:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd57;
                       end 
                      
                  9'd343/*343:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd56;
                       end 
                      
                  9'd344/*344:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd55;
                       end 
                      
                  9'd345/*345:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_ffff;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd54;
                       end 
                      
                  9'd346/*346:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd2;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd53;
                       end 
                      
                  9'd347/*347:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_ffff;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd52;
                       end 
                      
                  9'd348/*348:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd2;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd51;
                       end 
                      
                  9'd349/*349:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffd;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd50;
                       end 
                      
                  9'd350/*350:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffc;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd49;
                       end 
                      
                  9'd351/*351:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd48;
                       end 
                      
                  9'd352/*352:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd47;
                       end 
                      
                  9'd353/*353:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd1;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd46;
                       end 
                      
                  9'd354/*354:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd1;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd45;
                       end 
                      
                  9'd355/*355:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffa;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd44;
                       end 
                      
                  9'd356/*356:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd3;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd43;
                       end 
                      
                  9'd357/*357:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd4;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd42;
                       end 
                      
                  9'd358/*358:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffb;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd41;
                       end 
                      
                  9'd359/*359:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd40;
                       end 
                      
                  9'd360/*360:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd39;
                       end 
                      
                  9'd361/*361:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fff8;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd38;
                       end 
                      
                  9'd362/*362:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd37;
                       end 
                      
                  9'd363/*363:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd36;
                       end 
                      
                  9'd364/*364:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd35;
                       end 
                      
                  9'd365/*365:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffc;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd34;
                       end 
                      
                  9'd366/*366:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffb;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd33;
                       end 
                      
                  9'd367/*367:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffd;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd32;
                       end 
                      
                  9'd368/*368:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffc;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd31;
                       end 
                      
                  9'd369/*369:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffb;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd30;
                       end 
                      
                  9'd370/*370:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffa;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd29;
                       end 
                      
                  9'd371/*371:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffb;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd28;
                       end 
                      
                  9'd372/*372:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd27;
                       end 
                      
                  9'd373/*373:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffd;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd26;
                       end 
                      
                  9'd374/*374:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffd;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd25;
                       end 
                      
                  9'd375/*375:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffc;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd24;
                       end 
                      
                  9'd376/*376:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffb;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd23;
                       end 
                      
                  9'd377/*377:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffb;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd22;
                       end 
                      
                  9'd378/*378:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd12;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd21;
                       end 
                      
                  9'd379/*379:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd20;
                       end 
                      
                  9'd380/*380:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffd;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd19;
                       end 
                      
                  9'd381/*381:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_ffff;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd18;
                       end 
                      
                  9'd382/*382:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd17;
                       end 
                      
                  9'd383/*383:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd1;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd16;
                       end 
                      
                  9'd384/*384:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd1;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd15;
                       end 
                      
                  9'd385/*385:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd14;
                       end 
                      
                  9'd386/*386:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd13;
                       end 
                      
                  9'd387/*387:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd1;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd12;
                       end 
                      
                  9'd388/*388:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd11;
                       end 
                      
                  9'd389/*389:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_ffff;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd10;
                       end 
                      
                  9'd390/*390:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd9;
                       end 
                      
                  9'd391/*391:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_ffff;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd8;
                       end 
                      
                  9'd392/*392:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_ffff;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd7;
                       end 
                      
                  9'd393/*393:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_ffff;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd6;
                       end 
                      
                  9'd394/*394:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd1;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd5;
                       end 
                      
                  9'd395/*395:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffc;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd4;
                       end 
                      
                  9'd396/*396:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd3;
                       end 
                      
                  9'd397/*397:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd0;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd2;
                       end 
                      
                  9'd398/*398:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'h_ffff_fffe;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd1;
                       end 
                      
                  9'd399/*399:US*/:  begin 
                       A_SINT_CC_SCALbx16_ARA0_WRD0 = 32'd2;
                       A_SINT_CC_SCALbx16_ARA0_AD0 = 10'd0;
                       end 
                      
                  9'd402/*402:US*/:  begin 
                       iuMULTIPLIER10_DD = A_SINT_CC_SCALbx40_d2dim0;
                       iuMULTIPLIER10_NN = 64'hffffffffffffffff&TSPsw1_2_V_0;
                       iuMULTIPLIER12_DD = A_SINT_CC_SCALbx42_d2dim0;
                       iuMULTIPLIER12_NN = 64'hffffffffffffffff&TSPsw1_2_V_0;
                       iuMULTIPLIER14_DD = A_SINT_CC_SCALbx44_d2dim0;
                       iuMULTIPLIER14_NN = 64'hffffffffffffffff&TSPsw1_2_V_0;
                       end 
                      
                  9'd403/*403:US*/:  begin 
                       iuMULTIPLIER14_DD = A_SINT_CC_SCALbx46_d2dim0;
                       iuMULTIPLIER14_NN = 64'hffffffffffffffff&TSPsw1_2_V_0;
                       end 
                      
                  9'd405/*405:US*/:  begin 
                       A_64_SS_CC_SCALbx52_ARA0_WRD0 = 64'h_ffff_ffff_ffff_fff6;
                       A_64_SS_CC_SCALbx52_ARA0_AD0 = 64'd0+iuMULTIPLIER10_RR;
                       A_64_SS_CC_SCALbx54_ARB0_WRD0 = 64'd0;
                       A_64_SS_CC_SCALbx54_ARB0_AD0 = 64'd0+iuMULTIPLIER12_RR;
                       A_64_SS_CC_SCALbx56_ARC0_WRD0 = 64'd0;
                       A_64_SS_CC_SCALbx56_ARC0_AD0 = 64'd0+iuMULTIPLIER14_RR;
                       A_64_SS_CC_SCALbx58_ARD0_WRD0 = 64'd0;
                       A_64_SS_CC_SCALbx58_ARD0_AD0 = 64'd0+iuMULTIPLIER14_RR;
                       end 
                      
                  9'd407/*407:US*/:  begin 
                       A_64_SS_CC_SCALbx52_ARA0_WRD0 = 64'h_ffff_ffff_ffff_fff6;
                       A_64_SS_CC_SCALbx52_ARA0_AD0 = (64'hffffffffffffffff&TSPsw1_2_V_1)+64'd0*A_SINT_CC_SCALbx40_d2dim0;
                       A_64_SS_CC_SCALbx54_ARB0_WRD0 = 64'd0;
                       A_64_SS_CC_SCALbx54_ARB0_AD0 = (64'hffffffffffffffff&TSPsw1_2_V_1)+64'd0*A_SINT_CC_SCALbx42_d2dim0;
                       A_64_SS_CC_SCALbx56_ARC0_WRD0 = 64'd0;
                       A_64_SS_CC_SCALbx56_ARC0_AD0 = (64'hffffffffffffffff&TSPsw1_2_V_1)+64'd0*A_SINT_CC_SCALbx44_d2dim0;
                       A_64_SS_CC_SCALbx58_ARD0_WRD0 = 64'd0;
                       A_64_SS_CC_SCALbx58_ARD0_AD0 = (64'hffffffffffffffff&TSPsw1_2_V_1)+64'd0*A_SINT_CC_SCALbx46_d2dim0;
                       end 
                      
                  9'd409/*409:US*/:  begin 
                       A_16_SS_CC_SCALbx10_ARA0_AD0 = TSPru0_12_V_1;
                       A_16_SS_CC_SCALbx12_ARB0_AD0 = TSPen0_17_V_0;
                       end 
                      
                  9'd411/*411:US*/:  begin 
                       iuMULTIPLIER12_DD = A_SINT_CC_SCALbx40_d2dim0;
                       iuMULTIPLIER12_NN = 64'hffffffffffffffff&TSPne2_10_V_1;
                       iuMULTIPLIER14_DD = A_SINT_CC_SCALbx42_d2dim0;
                       iuMULTIPLIER14_NN = 64'hffffffffffffffff&TSPne2_10_V_1;
                       end 
                      endcase
              if ((xpc10nz==9'd413/*413:US*/))  A_64_SS_CC_SCALbx54_ARB0_AD0 = iuMULTIPLIER14_RR+(64'hffffffffffffffff&32'd1+TSPne2_10_V_3
                  );

                  
              case (xpc10nz)
                  9'd414/*414:US*/:  begin 
                       A_64_SS_CC_SCALbx52_ARA0_WRD0 = 64'h_ffff_ffff_ffff_fff6+A_64_SS_CC_SCALbx54_ARB0_RDD0;
                       A_64_SS_CC_SCALbx52_ARA0_AD0 = iuMULTIPLIER12_RR+(64'hffffffffffffffff&32'd1+TSPne2_10_V_3);
                       end 
                      
                  9'd416/*416:US*/:  begin 
                       iuMULTIPLIER14_DD = A_SINT_CC_SCALbx32_d2dim0;
                       iuMULTIPLIER14_NN = 64'hffffffffffffffff&TSPne2_10_V_4;
                       end 
                      endcase
              if ((xpc10nz==9'd418/*418:US*/))  A_SINT_CC_SCALbx16_ARA0_AD0 = (64'hffffffffffffffff&TSPne2_10_V_2)+iuMULTIPLIER14_RR;
                   end 
              if ((xpc10nz==9'd419/*419:US*/))  begin 
              if (((64'hffffffffffffffff&TSPne2_10_V_7+A_SINT_CC_SCALbx16_ARA0_RDD0)>=64'd0) && !xpc10_stall)  begin 
                       A_64_SS_CC_SCALbx54_ARB0_WRD0 = TSPne2_10_V_7+A_SINT_CC_SCALbx16_ARA0_RDD0;
                       A_64_SS_CC_SCALbx54_ARB0_AD0 = (64'hffffffffffffffff&32'd1+TSPne2_10_V_3)+(64'hffffffffffffffff&TSPne2_10_V_1)*
                      A_SINT_CC_SCALbx42_d2dim0;

                       end 
                      if (((64'hffffffffffffffff&TSPne2_10_V_7+A_SINT_CC_SCALbx16_ARA0_RDD0)<64'd0) && !xpc10_stall)  begin 
                       A_64_SS_CC_SCALbx54_ARB0_WRD0 = 64'd0;
                       A_64_SS_CC_SCALbx54_ARB0_AD0 = (64'hffffffffffffffff&32'd1+TSPne2_10_V_3)+(64'hffffffffffffffff&TSPne2_10_V_1)*
                      A_SINT_CC_SCALbx42_d2dim0;

                       end 
                       end 
              if (!xpc10_stall)  begin 
              if ((xpc10nz==9'd422/*422:US*/))  begin 
                       iuMULTIPLIER14_DD = A_SINT_CC_SCALbx42_d2dim0;
                       iuMULTIPLIER14_NN = 64'hffffffffffffffff&TSPne2_10_V_0;
                       end 
                      if ((xpc10nz==9'd424/*424:US*/))  A_64_SS_CC_SCALbx54_ARB0_AD0 = (64'hffffffffffffffff&TSPne2_10_V_3)+iuMULTIPLIER14_RR
                  ;

                  
              case (xpc10nz)
                  9'd426/*426:US*/:  begin 
                       iuMULTIPLIER12_DD = A_SINT_CC_SCALbx46_d2dim0;
                       iuMULTIPLIER12_NN = 64'hffffffffffffffff&TSPne2_10_V_0;
                       iuMULTIPLIER14_DD = A_SINT_CC_SCALbx44_d2dim0;
                       iuMULTIPLIER14_NN = 64'hffffffffffffffff&TSPne2_10_V_0;
                       end 
                      
                  9'd428/*428:US*/:  begin 
                       A_64_SS_CC_SCALbx56_ARC0_AD0 = (64'hffffffffffffffff&TSPne2_10_V_3)+iuMULTIPLIER14_RR;
                       A_64_SS_CC_SCALbx58_ARD0_AD0 = (64'hffffffffffffffff&TSPne2_10_V_3)+iuMULTIPLIER12_RR;
                       end 
                      
                  9'd430/*430:US*/:  begin 
                       iuMULTIPLIER12_DD = A_SINT_CC_SCALbx40_d2dim0;
                       iuMULTIPLIER12_NN = 64'hffffffffffffffff&TSPne2_10_V_1;
                       iuMULTIPLIER14_DD = A_SINT_CC_SCALbx44_d2dim0;
                       iuMULTIPLIER14_NN = 64'hffffffffffffffff&TSPne2_10_V_1;
                       end 
                      
                  9'd432/*432:US*/:  begin 
                       A_64_SS_CC_SCALbx52_ARA0_AD0 = (64'hffffffffffffffff&TSPne2_10_V_3)+iuMULTIPLIER12_RR;
                       A_64_SS_CC_SCALbx56_ARC0_AD0 = (64'hffffffffffffffff&TSPne2_10_V_3)+iuMULTIPLIER14_RR;
                       end 
                      endcase
               end 
              if ((xpc10nz==9'd433/*433:US*/))  begin 
              if (((64'hffffffffffffffff&64'h_ffff_ffff_ffff_fffe+A_64_SS_CC_SCALbx56_ARC0_RDD0)>=A_64_SS_CC_SCALbx52_ARA0_RDD0) && !xpc10_stall
              )  begin 
                       A_64_SS_CC_SCALbx58_ARD0_WRD0 = 64'h_ffff_ffff_ffff_fffe+A_64_SS_CC_SCALbx56_ARC0_RDD0;
                       A_64_SS_CC_SCALbx58_ARD0_AD0 = (64'hffffffffffffffff&32'd1+TSPne2_10_V_3)+(64'hffffffffffffffff&TSPne2_10_V_1)*
                      A_SINT_CC_SCALbx46_d2dim0;

                       end 
                      if (((64'hffffffffffffffff&64'h_ffff_ffff_ffff_fffe+A_64_SS_CC_SCALbx56_ARC0_RDD0)<A_64_SS_CC_SCALbx52_ARA0_RDD0
              ) && !xpc10_stall)  begin 
                       A_64_SS_CC_SCALbx56_ARC0_WRD0 = A_64_SS_CC_SCALbx52_ARA0_RDD0;
                       A_64_SS_CC_SCALbx56_ARC0_AD0 = iuMULTIPLIER14_RR+(64'hffffffffffffffff&32'd1+TSPne2_10_V_3);
                       end 
                       end 
              if (!xpc10_stall) 
          case (xpc10nz)
              9'd436/*436:US*/:  begin 
                   iuMULTIPLIER12_DD = A_SINT_CC_SCALbx40_d2dim0;
                   iuMULTIPLIER12_NN = 64'hffffffffffffffff&TSPne2_10_V_0;
                   iuMULTIPLIER14_DD = A_SINT_CC_SCALbx46_d2dim0;
                   iuMULTIPLIER14_NN = 64'hffffffffffffffff&TSPne2_10_V_0;
                   end 
                  
              9'd438/*438:US*/:  begin 
                   A_64_SS_CC_SCALbx52_ARA0_AD0 = iuMULTIPLIER12_RR+(64'hffffffffffffffff&32'd1+TSPne2_10_V_3);
                   A_64_SS_CC_SCALbx58_ARD0_AD0 = iuMULTIPLIER14_RR+(64'hffffffffffffffff&32'd1+TSPne2_10_V_3);
                   end 
                  endcase
          if ((xpc10nz==9'd439/*439:US*/))  begin 
              if (((64'hffffffffffffffff&64'h_ffff_ffff_ffff_fffe+A_64_SS_CC_SCALbx58_ARD0_RDD0)>=A_64_SS_CC_SCALbx52_ARA0_RDD0) && !xpc10_stall
              )  begin 
                       A_64_SS_CC_SCALbx58_ARD0_WRD0 = 64'h_ffff_ffff_ffff_fffe+A_64_SS_CC_SCALbx58_ARD0_RDD0;
                       A_64_SS_CC_SCALbx58_ARD0_AD0 = (64'hffffffffffffffff&32'd1+TSPne2_10_V_3)+(64'hffffffffffffffff&TSPne2_10_V_1)*
                      A_SINT_CC_SCALbx46_d2dim0;

                       end 
                      if (((64'hffffffffffffffff&64'h_ffff_ffff_ffff_fffe+A_64_SS_CC_SCALbx58_ARD0_RDD0)<A_64_SS_CC_SCALbx52_ARA0_RDD0
              ) && !xpc10_stall)  begin 
                       A_64_SS_CC_SCALbx58_ARD0_WRD0 = A_64_SS_CC_SCALbx52_ARA0_RDD0;
                       A_64_SS_CC_SCALbx58_ARD0_AD0 = (64'hffffffffffffffff&32'd1+TSPne2_10_V_3)+(64'hffffffffffffffff&TSPne2_10_V_1)*
                      A_SINT_CC_SCALbx46_d2dim0;

                       end 
                       end 
              if (!xpc10_stall)  begin 
              if ((xpc10nz==9'd442/*442:US*/))  begin 
                       iuMULTIPLIER14_DD = A_SINT_CC_SCALbx42_d2dim0;
                       iuMULTIPLIER14_NN = 64'hffffffffffffffff&TSPte2_13_V_1;
                       end 
                      if ((xpc10nz==9'd444/*444:US*/))  A_64_SS_CC_SCALbx54_ARB0_AD0 = (64'hffffffffffffffff&TSPte2_13_V_2)+iuMULTIPLIER14_RR
                  ;

                  if ((xpc10nz==9'd447/*447:US*/))  A_UINT_CC_SCALbx34_ARA0_AD0 = 8'hff&8'd255&32'hffffffff&TSPcr2_16_V_2;
                  if ((xpc10nz==9'd448/*448:US*/))  A_UINT_CC_SCALbx34_ARA0_AD0 = TCpr0_35_V_0;
                  if ((xpc10nz==9'd450/*450:US*/))  A_UINT_CC_SCALbx34_ARA0_AD0 = 8'hff&8'd255&((32'hffffffff&TSPcr2_16_V_2)>>5'd16);
                  if ((xpc10nz==9'd451/*451:US*/))  A_UINT_CC_SCALbx34_ARA0_AD0 = TCpr0_29_V_0;
                  if ((xpc10nz==9'd453/*453:US*/))  A_UINT_CC_SCALbx34_ARA0_AD0 = 8'hff&8'd255&((32'hffffffff&TSPcr2_16_V_2)>>4'd8);
                  if ((xpc10nz==9'd454/*454:US*/))  A_UINT_CC_SCALbx34_ARA0_AD0 = TCpr0_21_V_0;
                  if ((xpc10nz==9'd456/*456:US*/))  A_UINT_CC_SCALbx34_ARA0_AD0 = 8'hff&8'd255&32'hffffffff&TSPcr2_16_V_2;
                  if ((xpc10nz==9'd457/*457:US*/))  A_UINT_CC_SCALbx34_ARA0_AD0 = TCpr0_13_V_0;
                   end 
              if ((TSPcr2_16_V_1<32'd77) && !xpc10_stall)  begin 
              if ((xpc10nz==9'd459/*459:US*/))  begin 
                       iuMULTIPLIER14_DD = A_SINT_CC_SCALbx42_d2dim0;
                       iuMULTIPLIER14_NN = 64'hffffffffffffffff&TSPcr2_16_V_0;
                       end 
                      if ((xpc10nz==9'd461/*461:US*/))  A_64_SS_CC_SCALbx54_ARB0_AD0 = (64'hffffffffffffffff&TSPcr2_16_V_1)+iuMULTIPLIER14_RR
                  ;

                   end 
              if (!xpc10_stall)  begin 
              if ((xpc10nz==9'd473/*473:US*/))  A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd1;
                  if ((xpc10nz==9'd474/*474:US*/))  A_UINT_CC_SCALbx34_ARA0_AD0 = TCpr0_44_V_0;
                  if ((xpc10nz==9'd477/*477:US*/))  A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd128;
                  if ((xpc10nz==9'd478/*478:US*/))  A_UINT_CC_SCALbx34_ARA0_AD0 = TCpr0_40_V_0;
                  if ((xpc10nz==9'd481/*481:US*/))  A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd1;
                  if ((xpc10nz==9'd482/*482:US*/))  A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd255;
                  if ((xpc10nz==9'd484/*484:US*/))  A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd255;
                  if ((xpc10nz==9'd487/*487:US*/))  A_UINT_CC_SCALbx34_ARA0_AD0 = 9'd255;
                   end 
              if ((xpc10nz==9'd492/*492:US*/))  begin 
              if (((32'hffffffff&32'd1+TSPin0_6_V_0)<32'd77) && !xpc10_stall)  begin 
                       A_SINT_CC_SCALbx26_ARJ0_WRD0 = TSPe1_SPILL_256;
                       A_SINT_CC_SCALbx26_ARJ0_AD0 = TSPin0_6_V_0;
                       end 
                      if (((32'hffffffff&32'd1+TSPin0_6_V_0)>=32'd77) && !xpc10_stall)  begin 
                       A_SINT_CC_SCALbx26_ARJ0_WRD0 = TSPe1_SPILL_256;
                       A_SINT_CC_SCALbx26_ARJ0_AD0 = TSPin0_6_V_0;
                       end 
                       end 
              if ((xpc10nz==9'd495/*495:US*/) && !xpc10_stall)  begin 
               A_16_SS_CC_SCALbx14_ARC0_AD0 = TSPin0_6_V_0;
               A_16_SS_CC_SCALbx12_ARB0_AD0 = TSPen1_8_V_0;
               end 
               end 
      

 always   @(posedge clk )  begin 
      //Start structure HPR sw_test.exe
      if (reset)  begin 
               TCpr0_40_V_0 <= 8'd0;
               TCpr0_44_V_0 <= 8'd0;
               A_UINT_CC_SCALbx38_byteno <= 32'd0;
               A_UINT_CC_SCALbx38_crc_reg <= 32'd0;
               TSPru0_12_V_0 <= 32'd0;
               TSPne2_10_V_0 <= 32'd0;
               TSPne2_10_V_1 <= 32'd0;
               TSPne2_10_V_2 <= 32'd0;
               TSPte2_13_V_1 <= 32'd0;
               TSPcr2_16_V_0 <= 32'd0;
               TSPru0_12_V_1 <= 32'd0;
               TSPcr2_16_V_2 <= 64'd0;
               TCpr0_13_V_0 <= 8'd0;
               TCpr0_21_V_0 <= 8'd0;
               TCpr0_29_V_0 <= 8'd0;
               TCpr0_35_V_0 <= 8'd0;
               A_UINT_CC_SCALbx36_byteno <= 32'd0;
               A_UINT_CC_SCALbx36_crc_reg <= 32'd0;
               TSPcr2_16_V_1 <= 32'd0;
               TSPte2_13_V_0 <= 32'd0;
               TSPte2_13_V_2 <= 32'd0;
               TSPne2_10_V_4 <= 32'd0;
               TSPne2_10_V_7 <= 64'd0;
               TSPne2_10_V_3 <= 32'd0;
               TSPe0_SPILL_256 <= 32'd0;
               TSPen0_17_V_0 <= 32'd0;
               TSPsw1_2_V_1 <= 32'd0;
               d_monitor <= 64'd0;
               TSPsw1_2_V_0 <= 32'd0;
               TSPe1_SPILL_256 <= 32'd0;
               A_SINT_CC_SCALbx32_d2dim0 <= 32'd0;
               A_SINT_CC_SCALbx46_d2dim0 <= 32'd0;
               A_SINT_CC_SCALbx44_d2dim0 <= 32'd0;
               A_SINT_CC_SCALbx42_d2dim0 <= 32'd0;
               A_SINT_CC_SCALbx40_d2dim0 <= 32'd0;
               phase <= 32'd0;
               TSPin0_6_V_0 <= 32'd0;
               TSPen1_8_V_0 <= 32'd0;
               iuMULTIPLIER10RRh10hold <= 32'd0;
               iuMULTIPLIER10RRh10shot1 <= 1'd0;
               iuMULTIPLIER14RRh10hold <= 32'd0;
               iuMULTIPLIER14RRh10shot1 <= 1'd0;
               Z16SSCCSCALbx10ARA0RRh10hold <= 16'd0;
               SINTCCSCALbx16ARA0RRh10hold <= 32'd0;
               Z64SSCCSCALbx56ARC0RRh10hold <= 64'd0;
               iuMULTIPLIER12RRh10hold <= 32'd0;
               iuMULTIPLIER12RRh10shot1 <= 1'd0;
               Z64SSCCSCALbx52ARA0RRh10hold <= 64'd0;
               Z64SSCCSCALbx58ARD0RRh10hold <= 64'd0;
               iuMULTIPLIER14RRh12hold <= 32'd0;
               iuMULTIPLIER14RRh12shot1 <= 1'd0;
               Z64SSCCSCALbx54ARB0RRh10hold <= 64'd0;
               UINTCCSCALbx34ARA0RRh10hold <= 32'd0;
               UINTCCSCALbx34ARA0RRh12hold <= 32'd0;
               Z16SSCCSCALbx14ARC0RRh10hold <= 16'd0;
               Z16SSCCSCALbx12ARB0RRh10hold <= 16'd0;
               Z16SSCCSCALbx12ARB0RRh10shot0 <= 1'd0;
               Z16SSCCSCALbx14ARC0RRh10shot0 <= 1'd0;
               UINTCCSCALbx34ARA0RRh12shot0 <= 1'd0;
               UINTCCSCALbx34ARA0RRh10shot0 <= 1'd0;
               Z64SSCCSCALbx54ARB0RRh10shot0 <= 1'd0;
               iuMULTIPLIER14RRh12shot0 <= 1'd0;
               Z64SSCCSCALbx58ARD0RRh10shot0 <= 1'd0;
               Z64SSCCSCALbx52ARA0RRh10shot0 <= 1'd0;
               iuMULTIPLIER12RRh10shot0 <= 1'd0;
               Z64SSCCSCALbx56ARC0RRh10shot0 <= 1'd0;
               SINTCCSCALbx16ARA0RRh10shot0 <= 1'd0;
               Z16SSCCSCALbx10ARA0RRh10shot0 <= 1'd0;
               iuMULTIPLIER14RRh10shot0 <= 1'd0;
               iuMULTIPLIER10RRh10shot0 <= 1'd0;
               xpc10nz <= 9'd0;
               end 
               else  begin 
              if (((32'hffffffff&32'd1+TSPin0_6_V_0)>=32'd77) && (xpc10nz==9'd492/*492:US*/) && !xpc10_stall) $display("waypoint %1d %1d"
                  , 2'd3, 0);
                  if ((TSPru0_12_V_0>=32'd1) && (xpc10nz==9'd491/*491:US*/) && !xpc10_stall)  begin 
                      $display("waypoint %1d %1d", 4'd12, 0);
                      $display("CRC RESET");
                      $display("crc reg now:  reg=%H", 32'h_ffff_ffff);
                       end 
                      if (!xpc10_stall) 
                  case (xpc10nz)
                      9'd472/*472:US*/:  begin 
                          $display("self test yields %1d (should be 821105832)", A_UINT_CC_SCALbx38_crc_reg);
                          $display("Smith Waterman Simple Test End.");
                          $finish(0);
                           end 
                          
                      9'd475/*475:US*/:  begin 
                          $display("crc no=%1d dd=%1d cc=%H", A_UINT_CC_SCALbx38_byteno, 1'd1, TCpr0_44_V_0);
                          $display("crc update hex:  reg=%H,  tab[dd]=%H,  tab[cc]=%H", A_UINT_CC_SCALbx38_crc_reg, A_UINT_CC_SCALbx34_ARA0_RDD0
                          , A_UINT_CC_SCALbx34_ARA0_RDD0);
                           end 
                          
                      9'd479/*479:US*/:  begin 
                          $display("crc no=%1d dd=%1d cc=%H", A_UINT_CC_SCALbx38_byteno, 8'd128, TCpr0_40_V_0);
                          $display("crc update hex:  reg=%H,  tab[dd]=%H,  tab[cc]=%H", A_UINT_CC_SCALbx38_crc_reg, A_UINT_CC_SCALbx34_ARA0_RDD0
                          , A_UINT_CC_SCALbx34_ARA0_RDD0);
                           end 
                          
                      9'd483/*483:US*/:  begin 
                          $display("crc no=%1d dd=%1d cc=%H", A_UINT_CC_SCALbx38_byteno, 1'd1, 8'd255);
                          $display("crc update hex:  reg=%H,  tab[dd]=%H,  tab[cc]=%H", A_UINT_CC_SCALbx38_crc_reg, A_UINT_CC_SCALbx34_ARA0_RDD0
                          , A_UINT_CC_SCALbx34_ARA0_RDD0);
                           end 
                          
                      9'd485/*485:US*/: $display("self test startup %1d c ", A_UINT_CC_SCALbx34_ARA0_RDD0);

                      9'd486/*486:US*/: $display("self test startup %1d b ", 8'd255);

                      9'd488/*488:US*/: $display("self test startup %1d a ", A_UINT_CC_SCALbx34_ARA0_RDD0);
                  endcase
                  if ((TSPru0_12_V_1<2'd3) && (xpc10nz==9'd468/*468:US*/) && !xpc10_stall)  begin 
                      $display("waypoint %1d %1d", 3'd6, TSPru0_12_V_1);
                      $display("waypoint %1d %1d", 3'd4, 0);
                       end 
                      if ((TSPne2_10_V_3>=32'd77) && (xpc10nz==9'd465/*465:US*/) && !xpc10_stall)  begin 
                      $display("waypoint %1d %1d", 4'd8, TSPru0_12_V_1);
                      $display("Scored h matrix %1d", TSPru0_12_V_1);
                       end 
                      if ((TSPte2_13_V_0>=2'd2) && (xpc10nz==9'd464/*464:US*/) && !xpc10_stall)  begin 
                      $display("waypoint %1d %1d", 4'd10, TSPru0_12_V_1);
                      $display("CRC RESET");
                      $display("crc reg now:  reg=%H", 32'h_ffff_ffff);
                       end 
                      if ((TSPcr2_16_V_1>=32'd77) && (xpc10nz==9'd459/*459:US*/) && !xpc10_stall) $display("step %1d crc is %1d    0x%H"
                  , TSPru0_12_V_1, A_UINT_CC_SCALbx36_crc_reg, A_UINT_CC_SCALbx36_crc_reg);
                  if ((TSPcr2_16_V_1<32'd77) && (xpc10nz==9'd462/*462:US*/) && !xpc10_stall) $display("process unit word %1d word=%1d"
                  , A_UINT_CC_SCALbx36_byteno, 64'hffffffffffffffff&A_64_SS_CC_SCALbx54_ARB0_RDD0);
                  if (!xpc10_stall) 
                  case (xpc10nz)
                      0/*0:US*/:  begin 
                          $display("Smith Waterman Simple Test Start. Iterations=%1d", 32'd1);
                          $display("waypoint %1d %1d", 2'd2, 0);
                           A_SINT_CC_SCALbx32_d2dim0 <= 64'd20;
                           A_SINT_CC_SCALbx46_d2dim0 <= 32'd78;
                           A_SINT_CC_SCALbx44_d2dim0 <= 32'd78;
                           A_SINT_CC_SCALbx42_d2dim0 <= 32'd78;
                           A_SINT_CC_SCALbx40_d2dim0 <= 32'd78;
                           phase <= 32'd2;
                           TSPin0_6_V_0 <= 32'd0;
                           TSPen1_8_V_0 <= 32'd0;
                           end 
                          
                      9'd405/*405:US*/:  begin 
                           d_monitor <= TSPsw1_2_V_0;
                           TSPsw1_2_V_0 <= 32'd1+TSPsw1_2_V_0;
                           end 
                          
                      9'd407/*407:US*/:  TSPsw1_2_V_1 <= 32'd1+TSPsw1_2_V_1;

                      9'd414/*414:US*/:  TSPne2_10_V_3 <= 32'd1+TSPne2_10_V_3;

                      9'd445/*445:US*/:  begin 
                          $write("%1d %1d : %1d   ", TSPte2_13_V_1, TSPte2_13_V_2, 64'hffffffffffffffff&A_64_SS_CC_SCALbx54_ARB0_RDD0
                          );
                          $display("");
                           TSPte2_13_V_2 <= 32'd1+TSPte2_13_V_2;
                           end 
                          
                      9'd449/*449:US*/:  begin 
                          $display("crc no=%1d dd=%1d cc=%H", A_UINT_CC_SCALbx36_byteno, 8'hff&8'd255&32'hffffffff&TSPcr2_16_V_2, TCpr0_35_V_0
                          );
                          $display("crc update hex:  reg=%H,  tab[dd]=%H,  tab[cc]=%H", A_UINT_CC_SCALbx36_crc_reg, A_UINT_CC_SCALbx34_ARA0_RDD0
                          , A_UINT_CC_SCALbx34_ARA0_RDD0);
                           A_UINT_CC_SCALbx36_crc_reg <= -32'd1&{A_UINT_CC_SCALbx36_crc_reg, 8'd0};
                           TSPcr2_16_V_1 <= 32'd1+TSPcr2_16_V_1;
                           end 
                          
                      9'd452/*452:US*/:  begin 
                          $display("crc no=%1d dd=%1d cc=%H", A_UINT_CC_SCALbx36_byteno, 8'hff&8'd255&((32'hffffffff&TSPcr2_16_V_2)>>
                          5'd16), TCpr0_29_V_0);
                          $display("crc update hex:  reg=%H,  tab[dd]=%H,  tab[cc]=%H", A_UINT_CC_SCALbx36_crc_reg, A_UINT_CC_SCALbx34_ARA0_RDD0
                          , A_UINT_CC_SCALbx34_ARA0_RDD0);
                           TCpr0_35_V_0 <= 8'd255&((32'hffffffff&-32'd1&{A_UINT_CC_SCALbx36_crc_reg, 8'd0})>>5'd24);
                           A_UINT_CC_SCALbx36_byteno <= 32'd1+A_UINT_CC_SCALbx36_byteno;
                           A_UINT_CC_SCALbx36_crc_reg <= -32'd1&{A_UINT_CC_SCALbx36_crc_reg, 8'd0};
                           end 
                          
                      9'd455/*455:US*/:  begin 
                          $display("crc no=%1d dd=%1d cc=%H", A_UINT_CC_SCALbx36_byteno, 8'hff&8'd255&((32'hffffffff&TSPcr2_16_V_2)>>
                          4'd8), TCpr0_21_V_0);
                          $display("crc update hex:  reg=%H,  tab[dd]=%H,  tab[cc]=%H", A_UINT_CC_SCALbx36_crc_reg, A_UINT_CC_SCALbx34_ARA0_RDD0
                          , A_UINT_CC_SCALbx34_ARA0_RDD0);
                           TCpr0_29_V_0 <= 8'd255&((32'hffffffff&-32'd1&{A_UINT_CC_SCALbx36_crc_reg, 8'd0})>>5'd24);
                           A_UINT_CC_SCALbx36_byteno <= 32'd1+A_UINT_CC_SCALbx36_byteno;
                           A_UINT_CC_SCALbx36_crc_reg <= -32'd1&{A_UINT_CC_SCALbx36_crc_reg, 8'd0};
                           end 
                          
                      9'd458/*458:US*/:  begin 
                          $display("crc no=%1d dd=%1d cc=%H", A_UINT_CC_SCALbx36_byteno, 8'hff&8'd255&32'hffffffff&TSPcr2_16_V_2, TCpr0_13_V_0
                          );
                          $display("crc update hex:  reg=%H,  tab[dd]=%H,  tab[cc]=%H", A_UINT_CC_SCALbx36_crc_reg, A_UINT_CC_SCALbx34_ARA0_RDD0
                          , A_UINT_CC_SCALbx34_ARA0_RDD0);
                           TCpr0_21_V_0 <= 8'd255&((32'hffffffff&-32'd1&{A_UINT_CC_SCALbx36_crc_reg, 8'd0})>>5'd24);
                           A_UINT_CC_SCALbx36_byteno <= 32'd1+A_UINT_CC_SCALbx36_byteno;
                           A_UINT_CC_SCALbx36_crc_reg <= -32'd1&{A_UINT_CC_SCALbx36_crc_reg, 8'd0};
                           end 
                          
                      9'd463/*463:US*/:  begin 
                           TSPcr2_16_V_0 <= ((32'd1+TSPru0_12_V_1)%2'd2);
                           TSPcr2_16_V_1 <= 32'd0;
                           end 
                          
                      9'd466/*466:US*/:  begin 
                           TSPne2_10_V_2 <= TSPe0_SPILL_256;
                           TSPne2_10_V_3 <= 32'd0;
                           end 
                          
                      9'd471/*471:US*/:  TSPsw1_2_V_0 <= 32'd0;

                      9'd475/*475:US*/:  A_UINT_CC_SCALbx38_crc_reg <= -32'd1&{A_UINT_CC_SCALbx38_crc_reg, 8'd0};

                      9'd476/*476:US*/:  begin 
                           TCpr0_44_V_0 <= 8'd255&(A_UINT_CC_SCALbx38_crc_reg>>5'd24);
                           A_UINT_CC_SCALbx38_byteno <= 32'd1+A_UINT_CC_SCALbx38_byteno;
                           end 
                          
                      9'd479/*479:US*/:  A_UINT_CC_SCALbx38_crc_reg <= -32'd1&{A_UINT_CC_SCALbx38_crc_reg, 8'd0};

                      9'd480/*480:US*/:  begin 
                           TCpr0_40_V_0 <= 8'd255&(A_UINT_CC_SCALbx38_crc_reg>>5'd24);
                           A_UINT_CC_SCALbx38_byteno <= 32'd1+A_UINT_CC_SCALbx38_byteno;
                           end 
                          
                      9'd483/*483:US*/:  A_UINT_CC_SCALbx38_crc_reg <= -32'd1&{A_UINT_CC_SCALbx38_crc_reg, 8'd0};

                      9'd485/*485:US*/:  A_UINT_CC_SCALbx38_byteno <= 32'd1+A_UINT_CC_SCALbx38_byteno;

                      9'd489/*489:US*/:  A_UINT_CC_SCALbx38_crc_reg <= 32'h_ffff_ffff;
                  endcase
                  if (UINTCCSCALbx34ARA0RRh12shot0)  begin 
                      
                      case (xpc10nz)
                          9'd449/*449:US*/:  xpc10nz <= 9'd459/*459:xpc10nz*/;

                          9'd485/*485:US*/:  xpc10nz <= 9'd481/*481:xpc10nz*/;

                          9'd488/*488:US*/:  xpc10nz <= 9'd486/*486:xpc10nz*/;
                      endcase
                       UINTCCSCALbx34ARA0RRh12hold <= A_UINT_CC_SCALbx34_ARA0_RDD0;
                       UINTCCSCALbx34ARA0RRh12hold <= A_UINT_CC_SCALbx34_ARA0_RDD0;
                       UINTCCSCALbx34ARA0RRh12hold <= A_UINT_CC_SCALbx34_ARA0_RDD0;
                       UINTCCSCALbx34ARA0RRh12hold <= A_UINT_CC_SCALbx34_ARA0_RDD0;
                       UINTCCSCALbx34ARA0RRh12hold <= A_UINT_CC_SCALbx34_ARA0_RDD0;
                       UINTCCSCALbx34ARA0RRh12hold <= A_UINT_CC_SCALbx34_ARA0_RDD0;
                       UINTCCSCALbx34ARA0RRh12hold <= A_UINT_CC_SCALbx34_ARA0_RDD0;
                      if ((xpc10nz==9'd451/*451:US*/))  xpc10nz <= 9'd452/*452:xpc10nz*/;
                          if ((xpc10nz==9'd454/*454:US*/))  xpc10nz <= 9'd455/*455:xpc10nz*/;
                          if ((xpc10nz==9'd457/*457:US*/))  xpc10nz <= 9'd458/*458:xpc10nz*/;
                          if ((xpc10nz==9'd474/*474:US*/))  xpc10nz <= 9'd475/*475:xpc10nz*/;
                          if ((xpc10nz==9'd478/*478:US*/))  xpc10nz <= 9'd479/*479:xpc10nz*/;
                          if ((xpc10nz==9'd482/*482:US*/))  xpc10nz <= 9'd483/*483:xpc10nz*/;
                           end 
                      if (UINTCCSCALbx34ARA0RRh10shot0)  begin 
                      
                      case (xpc10nz)
                          9'd452/*452:US*/:  xpc10nz <= 9'd447/*447:xpc10nz*/;

                          9'd455/*455:US*/:  xpc10nz <= 9'd450/*450:xpc10nz*/;

                          9'd458/*458:US*/:  xpc10nz <= 9'd453/*453:xpc10nz*/;

                          9'd475/*475:US*/:  xpc10nz <= 9'd472/*472:xpc10nz*/;

                          9'd479/*479:US*/:  xpc10nz <= 9'd476/*476:xpc10nz*/;

                          9'd483/*483:US*/:  xpc10nz <= 9'd480/*480:xpc10nz*/;
                      endcase
                       UINTCCSCALbx34ARA0RRh10hold <= A_UINT_CC_SCALbx34_ARA0_RDD0;
                       UINTCCSCALbx34ARA0RRh10hold <= A_UINT_CC_SCALbx34_ARA0_RDD0;
                       UINTCCSCALbx34ARA0RRh10hold <= A_UINT_CC_SCALbx34_ARA0_RDD0;
                       UINTCCSCALbx34ARA0RRh10hold <= A_UINT_CC_SCALbx34_ARA0_RDD0;
                       UINTCCSCALbx34ARA0RRh10hold <= A_UINT_CC_SCALbx34_ARA0_RDD0;
                       UINTCCSCALbx34ARA0RRh10hold <= A_UINT_CC_SCALbx34_ARA0_RDD0;
                       UINTCCSCALbx34ARA0RRh10hold <= A_UINT_CC_SCALbx34_ARA0_RDD0;
                      if ((xpc10nz==9'd448/*448:US*/))  xpc10nz <= 9'd449/*449:xpc10nz*/;
                           end 
                      if ((xpc10nz==0/*0:US*/))  xpc10nz <= 1'd1/*1:xpc10nz*/;
                  if (iuMULTIPLIER14RRh12shot1)  begin 
                       iuMULTIPLIER14RRh12hold <= iuMULTIPLIER14_RR;
                       iuMULTIPLIER14RRh12hold <= iuMULTIPLIER14_RR;
                       iuMULTIPLIER14RRh12hold <= iuMULTIPLIER14_RR;
                       iuMULTIPLIER14RRh12hold <= iuMULTIPLIER14_RR;
                       iuMULTIPLIER14RRh12hold <= iuMULTIPLIER14_RR;
                       iuMULTIPLIER14RRh12hold <= iuMULTIPLIER14_RR;
                       iuMULTIPLIER14RRh12hold <= iuMULTIPLIER14_RR;
                       iuMULTIPLIER14RRh12hold <= iuMULTIPLIER14_RR;
                       iuMULTIPLIER14RRh12hold <= iuMULTIPLIER14_RR;
                       end 
                      
              case (xpc10nz)
                  9'd464/*464:US*/:  begin 
                      if ((TSPte2_13_V_0>=2'd2) && !xpc10_stall)  begin 
                               A_UINT_CC_SCALbx36_crc_reg <= 32'h_ffff_ffff;
                               phase <= 32'd10+32'd256*TSPru0_12_V_1;
                               end 
                              if ((TSPte2_13_V_0<2'd2))  xpc10nz <= 9'd446/*446:xpc10nz*/;
                           else  xpc10nz <= 9'd463/*463:xpc10nz*/;
                      if ((TSPte2_13_V_0<2'd2) && !xpc10_stall)  begin 
                               TSPte2_13_V_1 <= ((TSPru0_12_V_1+TSPte2_13_V_0)%2'd2);
                               TSPte2_13_V_2 <= 32'd0;
                               end 
                               end 
                      
                  9'd468/*468:US*/:  begin 
                      if ((TSPru0_12_V_1<2'd3) && !xpc10_stall)  begin 
                               TSPne2_10_V_0 <= (TSPru0_12_V_1%2'd2);
                               TSPne2_10_V_1 <= ((32'd1+TSPru0_12_V_1)%2'd2);
                               TSPen0_17_V_0 <= 32'd0;
                               phase <= 32'd4;
                               end 
                              if ((TSPru0_12_V_1<2'd3))  xpc10nz <= 9'd467/*467:xpc10nz*/;
                           else  xpc10nz <= 9'd491/*491:xpc10nz*/;
                      if ((TSPru0_12_V_1>=2'd3) && !xpc10_stall)  TSPru0_12_V_0 <= 32'd1+TSPru0_12_V_0;
                           end 
                      endcase
              if (Z64SSCCSCALbx54ARB0RRh10shot0)  begin 
                      
                      case (xpc10nz)
                          9'd414/*414:US*/:  xpc10nz <= 9'd415/*415:xpc10nz*/;

                          9'd425/*425:US*/:  xpc10nz <= 9'd416/*416:xpc10nz*/;

                          9'd445/*445:US*/:  xpc10nz <= 9'd446/*446:xpc10nz*/;

                          9'd462/*462:US*/:  xpc10nz <= 9'd456/*456:xpc10nz*/;
                      endcase
                       Z64SSCCSCALbx54ARB0RRh10hold <= A_64_SS_CC_SCALbx54_ARB0_RDD0;
                       Z64SSCCSCALbx54ARB0RRh10hold <= A_64_SS_CC_SCALbx54_ARB0_RDD0;
                       Z64SSCCSCALbx54ARB0RRh10hold <= A_64_SS_CC_SCALbx54_ARB0_RDD0;
                       Z64SSCCSCALbx54ARB0RRh10hold <= A_64_SS_CC_SCALbx54_ARB0_RDD0;
                       end 
                      
              case (xpc10nz)
                  9'd465/*465:US*/:  begin 
                      if ((TSPne2_10_V_3>=32'd77) && !xpc10_stall)  begin 
                               TSPte2_13_V_0 <= 32'd0;
                               phase <= 32'd8+32'd256*TSPru0_12_V_1;
                               end 
                              if ((TSPne2_10_V_3<32'd77))  xpc10nz <= 9'd436/*436:xpc10nz*/;
                           else  xpc10nz <= 9'd464/*464:xpc10nz*/;
                       end 
                      
                  9'd491/*491:US*/:  begin 
                      if ((TSPru0_12_V_0>=32'd1) && !xpc10_stall)  begin 
                               A_UINT_CC_SCALbx38_crc_reg <= 32'h_ffff_ffff;
                               phase <= 32'd12;
                               end 
                              if ((TSPru0_12_V_0<32'd1))  xpc10nz <= 9'd471/*471:xpc10nz*/;
                           else  xpc10nz <= 9'd490/*490:xpc10nz*/;
                       end 
                      
                  9'd492/*492:US*/:  begin 
                      if (((32'hffffffff&32'd1+TSPin0_6_V_0)>=32'd77) && !xpc10_stall)  begin 
                               TSPru0_12_V_0 <= 32'd0;
                               phase <= 32'd3;
                               TSPin0_6_V_0 <= 32'd1+TSPin0_6_V_0;
                               end 
                              if (((32'hffffffff&32'd1+TSPin0_6_V_0)<32'd77))  xpc10nz <= 9'd494/*494:xpc10nz*/;
                           else  xpc10nz <= 9'd493/*493:xpc10nz*/;
                      if (((32'hffffffff&32'd1+TSPin0_6_V_0)<32'd77) && !xpc10_stall)  begin 
                               TSPin0_6_V_0 <= 32'd1+TSPin0_6_V_0;
                               TSPen1_8_V_0 <= 32'd0;
                               end 
                               end 
                      endcase
              if (iuMULTIPLIER12RRh10shot1)  begin 
                       iuMULTIPLIER12RRh10hold <= iuMULTIPLIER12_RR;
                       iuMULTIPLIER12RRh10hold <= iuMULTIPLIER12_RR;
                       iuMULTIPLIER12RRh10hold <= iuMULTIPLIER12_RR;
                       iuMULTIPLIER12RRh10hold <= iuMULTIPLIER12_RR;
                       iuMULTIPLIER12RRh10hold <= iuMULTIPLIER12_RR;
                       end 
                      if ((TSPcr2_16_V_1<32'd77) && (xpc10nz==9'd462/*462:US*/) && !xpc10_stall)  begin 
                       TSPcr2_16_V_2 <= A_64_SS_CC_SCALbx54_ARB0_RDD0;
                       TCpr0_13_V_0 <= 8'd255&(A_UINT_CC_SCALbx36_crc_reg>>5'd24);
                       A_UINT_CC_SCALbx36_byteno <= 32'd1+A_UINT_CC_SCALbx36_byteno;
                       end 
                      
              case (xpc10nz)
                  9'd401/*401:US*/:  begin 
                      if ((TSPen1_8_V_0<5'd20))  xpc10nz <= 9'd497/*497:xpc10nz*/;
                           else  xpc10nz <= 9'd492/*492:xpc10nz*/;
                      if ((TSPen1_8_V_0>=5'd20) && !xpc10_stall)  TSPe1_SPILL_256 <= 32'd0;
                           end 
                      
                  9'd405/*405:US*/:  xpc10nz <= 9'd406/*406:xpc10nz*/;

                  9'd410/*410:US*/:  begin 
                      if ((A_16_SS_CC_SCALbx10_ARA0_RDD0==A_16_SS_CC_SCALbx12_ARB0_RDD0) && !xpc10_stall)  TSPe0_SPILL_256 <= TSPen0_17_V_0
                          ;

                          if ((A_16_SS_CC_SCALbx10_ARA0_RDD0!=A_16_SS_CC_SCALbx12_ARB0_RDD0) && !xpc10_stall)  TSPen0_17_V_0 <= 32'd1
                          +TSPen0_17_V_0;

                          if (Z16SSCCSCALbx10ARA0RRh10shot0 && Z16SSCCSCALbx12ARB0RRh10shot0 && (A_16_SS_CC_SCALbx10_ARA0_RDD0==A_16_SS_CC_SCALbx12_ARB0_RDD0
                      ))  xpc10nz <= 9'd466/*466:xpc10nz*/;
                          if (Z16SSCCSCALbx10ARA0RRh10shot0 && Z16SSCCSCALbx12ARB0RRh10shot0 && (A_16_SS_CC_SCALbx10_ARA0_RDD0!=A_16_SS_CC_SCALbx12_ARB0_RDD0
                      ))  xpc10nz <= 9'd467/*467:xpc10nz*/;
                           end 
                      
                  9'd419/*419:US*/:  begin 
                      if (SINTCCSCALbx16ARA0RRh10shot0 && ((64'hffffffffffffffff&TSPne2_10_V_7+A_SINT_CC_SCALbx16_ARA0_RDD0)<64'd0)) 
                       xpc10nz <= 9'd420/*420:xpc10nz*/;
                          if (SINTCCSCALbx16ARA0RRh10shot0 && ((64'hffffffffffffffff&TSPne2_10_V_7+A_SINT_CC_SCALbx16_ARA0_RDD0)>=64'd0
                      ))  xpc10nz <= 9'd421/*421:xpc10nz*/;
                           end 
                      
                  9'd429/*429:US*/:  begin 
                      if ((A_64_SS_CC_SCALbx56_ARC0_RDD0<A_64_SS_CC_SCALbx58_ARD0_RDD0) && !xpc10_stall)  TSPne2_10_V_7 <= A_64_SS_CC_SCALbx58_ARD0_RDD0
                          ;

                          if ((A_64_SS_CC_SCALbx56_ARC0_RDD0>=A_64_SS_CC_SCALbx58_ARD0_RDD0) && !xpc10_stall)  TSPne2_10_V_7 <= A_64_SS_CC_SCALbx56_ARC0_RDD0
                          ;

                          if (Z64SSCCSCALbx56ARC0RRh10shot0 && Z64SSCCSCALbx58ARD0RRh10shot0)  xpc10nz <= 9'd422/*422:xpc10nz*/;
                           end 
                      
                  9'd433/*433:US*/:  begin 
                      if (Z64SSCCSCALbx56ARC0RRh10shot0 && Z64SSCCSCALbx52ARA0RRh10shot0 && ((64'hffffffffffffffff&64'h_ffff_ffff_ffff_fffe
                      +A_64_SS_CC_SCALbx56_ARC0_RDD0)<A_64_SS_CC_SCALbx52_ARA0_RDD0))  xpc10nz <= 9'd434/*434:xpc10nz*/;
                          if (Z64SSCCSCALbx56ARC0RRh10shot0 && Z64SSCCSCALbx52ARA0RRh10shot0 && ((64'hffffffffffffffff&64'h_ffff_ffff_ffff_fffe
                      +A_64_SS_CC_SCALbx56_ARC0_RDD0)>=A_64_SS_CC_SCALbx52_ARA0_RDD0))  xpc10nz <= 9'd435/*435:xpc10nz*/;
                           end 
                      
                  9'd439/*439:US*/:  begin 
                      if (((64'hffffffffffffffff&64'h_ffff_ffff_ffff_fffe+A_64_SS_CC_SCALbx58_ARD0_RDD0)<A_64_SS_CC_SCALbx52_ARA0_RDD0
                      ) && !xpc10_stall)  TSPne2_10_V_4 <= A_SINT_CC_SCALbx26_ARJ0[TSPne2_10_V_3];
                      if (((64'hffffffffffffffff&64'h_ffff_ffff_ffff_fffe+A_64_SS_CC_SCALbx58_ARD0_RDD0)>=A_64_SS_CC_SCALbx52_ARA0_RDD0
                      ) && !xpc10_stall)  TSPne2_10_V_4 <= A_SINT_CC_SCALbx26_ARJ0[TSPne2_10_V_3];

                          if (Z64SSCCSCALbx58ARD0RRh10shot0 && Z64SSCCSCALbx52ARA0RRh10shot0 && ((64'hffffffffffffffff&64'h_ffff_ffff_ffff_fffe
                      +A_64_SS_CC_SCALbx58_ARD0_RDD0)<A_64_SS_CC_SCALbx52_ARA0_RDD0))  xpc10nz <= 9'd440/*440:xpc10nz*/;
                          if (Z64SSCCSCALbx58ARD0RRh10shot0 && Z64SSCCSCALbx52ARA0RRh10shot0 && ((64'hffffffffffffffff&64'h_ffff_ffff_ffff_fffe
                      +A_64_SS_CC_SCALbx58_ARD0_RDD0)>=A_64_SS_CC_SCALbx52_ARA0_RDD0))  xpc10nz <= 9'd441/*441:xpc10nz*/;
                           end 
                      
                  9'd446/*446:US*/:  begin 
                      if ((TSPte2_13_V_2<32'd77))  xpc10nz <= 9'd442/*442:xpc10nz*/;
                           else  xpc10nz <= 9'd464/*464:xpc10nz*/;
                      if ((TSPte2_13_V_2>=32'd77) && !xpc10_stall)  TSPte2_13_V_0 <= 32'd1+TSPte2_13_V_0;
                           end 
                      
                  9'd459/*459:US*/:  begin 
                      if ((TSPcr2_16_V_1>=32'd77) && !xpc10_stall)  begin 
                               TSPru0_12_V_1 <= 32'd1+TSPru0_12_V_1;
                               d_monitor <= A_UINT_CC_SCALbx36_crc_reg;
                               end 
                              if ((TSPcr2_16_V_1<32'd77))  xpc10nz <= 9'd460/*460:xpc10nz*/;
                           else  xpc10nz <= 9'd468/*468:xpc10nz*/;
                       end 
                      
                  9'd463/*463:US*/:  xpc10nz <= 9'd459/*459:xpc10nz*/;

                  9'd466/*466:US*/:  xpc10nz <= 9'd465/*465:xpc10nz*/;

                  9'd467/*467:US*/:  begin 
                      if ((TSPen0_17_V_0<5'd20))  xpc10nz <= 9'd409/*409:xpc10nz*/;
                           else  xpc10nz <= 9'd466/*466:xpc10nz*/;
                      if ((TSPen0_17_V_0>=5'd20) && !xpc10_stall)  TSPe0_SPILL_256 <= 32'd0;
                           end 
                      
                  9'd469/*469:US*/:  begin 
                      if ((TSPsw1_2_V_1<7'd78))  xpc10nz <= 9'd407/*407:xpc10nz*/;
                           else  xpc10nz <= 9'd468/*468:xpc10nz*/;
                      if ((TSPsw1_2_V_1>=7'd78) && !xpc10_stall)  TSPru0_12_V_1 <= 32'd0;
                           end 
                      
                  9'd470/*470:US*/:  begin 
                      if ((TSPsw1_2_V_0<2'd2))  xpc10nz <= 9'd402/*402:xpc10nz*/;
                           else  xpc10nz <= 9'd469/*469:xpc10nz*/;
                      if ((TSPsw1_2_V_0>=2'd2) && !xpc10_stall)  TSPsw1_2_V_1 <= 32'd1;
                           end 
                      
                  9'd472/*472:US*/:  xpc10nz <= 9'd472/*472:xpc10nz*/;

                  9'd476/*476:US*/:  xpc10nz <= 9'd473/*473:xpc10nz*/;

                  9'd480/*480:US*/:  xpc10nz <= 9'd477/*477:xpc10nz*/;

                  9'd486/*486:US*/:  xpc10nz <= 9'd484/*484:xpc10nz*/;

                  9'd496/*496:US*/:  begin 
                      if ((A_16_SS_CC_SCALbx12_ARB0_RDD0==A_16_SS_CC_SCALbx14_ARC0_RDD0) && !xpc10_stall)  TSPe1_SPILL_256 <= TSPen1_8_V_0
                          ;

                          if ((A_16_SS_CC_SCALbx12_ARB0_RDD0!=A_16_SS_CC_SCALbx14_ARC0_RDD0) && !xpc10_stall)  TSPen1_8_V_0 <= 32'd1+
                          TSPen1_8_V_0;

                          if (Z16SSCCSCALbx12ARB0RRh10shot0 && Z16SSCCSCALbx14ARC0RRh10shot0 && (A_16_SS_CC_SCALbx12_ARB0_RDD0==A_16_SS_CC_SCALbx14_ARC0_RDD0
                      ))  xpc10nz <= 9'd492/*492:xpc10nz*/;
                          if (Z16SSCCSCALbx12ARB0RRh10shot0 && Z16SSCCSCALbx14ARC0RRh10shot0 && (A_16_SS_CC_SCALbx12_ARB0_RDD0!=A_16_SS_CC_SCALbx14_ARC0_RDD0
                      ))  xpc10nz <= 9'd401/*401:xpc10nz*/;
                           end 
                      endcase
              if (Z64SSCCSCALbx52ARA0RRh10shot0)  begin 
                       Z64SSCCSCALbx52ARA0RRh10hold <= A_64_SS_CC_SCALbx52_ARA0_RDD0;
                       Z64SSCCSCALbx52ARA0RRh10hold <= A_64_SS_CC_SCALbx52_ARA0_RDD0;
                       end 
                      if (Z64SSCCSCALbx58ARD0RRh10shot0)  begin 
                       Z64SSCCSCALbx58ARD0RRh10hold <= A_64_SS_CC_SCALbx58_ARD0_RDD0;
                       Z64SSCCSCALbx58ARD0RRh10hold <= A_64_SS_CC_SCALbx58_ARD0_RDD0;
                       end 
                      if (Z64SSCCSCALbx56ARC0RRh10shot0)  begin 
                       Z64SSCCSCALbx56ARC0RRh10hold <= A_64_SS_CC_SCALbx56_ARC0_RDD0;
                       Z64SSCCSCALbx56ARC0RRh10hold <= A_64_SS_CC_SCALbx56_ARC0_RDD0;
                       end 
                      if (Z16SSCCSCALbx12ARB0RRh10shot0)  begin 
                       Z16SSCCSCALbx12ARB0RRh10hold <= A_16_SS_CC_SCALbx12_ARB0_RDD0;
                       Z16SSCCSCALbx12ARB0RRh10hold <= A_16_SS_CC_SCALbx12_ARB0_RDD0;
                       end 
                      
              case (xpc10nz)
                  9'd407/*407:US*/:  xpc10nz <= 9'd408/*408:xpc10nz*/;

                  9'd425/*425:US*/: if ((TSPne2_10_V_7<A_64_SS_CC_SCALbx54_ARB0_RDD0) && !xpc10_stall)  TSPne2_10_V_7 <= A_64_SS_CC_SCALbx54_ARB0_RDD0
                      ;

                      
                  9'd471/*471:US*/:  xpc10nz <= 9'd470/*470:xpc10nz*/;

                  9'd489/*489:US*/:  xpc10nz <= 9'd487/*487:xpc10nz*/;
              endcase
              if (iuMULTIPLIER10RRh10shot1)  iuMULTIPLIER10RRh10hold <= iuMULTIPLIER10_RR;
                   iuMULTIPLIER10RRh10shot1 <= iuMULTIPLIER10RRh10shot0;
              if (iuMULTIPLIER14RRh10shot1)  iuMULTIPLIER14RRh10hold <= iuMULTIPLIER14_RR;
                   iuMULTIPLIER14RRh10shot1 <= iuMULTIPLIER14RRh10shot0;
              if (Z16SSCCSCALbx10ARA0RRh10shot0)  Z16SSCCSCALbx10ARA0RRh10hold <= A_16_SS_CC_SCALbx10_ARA0_RDD0;
                  if (SINTCCSCALbx16ARA0RRh10shot0)  SINTCCSCALbx16ARA0RRh10hold <= A_SINT_CC_SCALbx16_ARA0_RDD0;
                   iuMULTIPLIER12RRh10shot1 <= iuMULTIPLIER12RRh10shot0;
               iuMULTIPLIER14RRh12shot1 <= iuMULTIPLIER14RRh12shot0;
              if (Z16SSCCSCALbx14ARC0RRh10shot0)  Z16SSCCSCALbx14ARC0RRh10hold <= A_16_SS_CC_SCALbx14_ARC0_RDD0;
                   Z16SSCCSCALbx12ARB0RRh10shot0 <= ((xpc10nz==9'd495/*495:US*/) || (xpc10nz==9'd409/*409:US*/)) && !xpc10_stall;
               Z16SSCCSCALbx14ARC0RRh10shot0 <= (xpc10nz==9'd495/*495:US*/) && !xpc10_stall;
               UINTCCSCALbx34ARA0RRh12shot0 <= ((xpc10nz==9'd487/*487:US*/) || (xpc10nz==9'd481/*481:US*/) || (xpc10nz==9'd473/*473:US*/) || 
              (xpc10nz==9'd453/*453:US*/) || (xpc10nz==9'd448/*448:US*/) || (xpc10nz==9'd450/*450:US*/) || (xpc10nz==9'd456/*456:US*/) || 
              (xpc10nz==9'd477/*477:US*/) || (xpc10nz==9'd484/*484:US*/)) && !xpc10_stall;

               UINTCCSCALbx34ARA0RRh10shot0 <= ((xpc10nz==9'd482/*482:US*/) || (xpc10nz==9'd474/*474:US*/) || (xpc10nz==9'd454/*454:US*/) || 
              (xpc10nz==9'd447/*447:US*/) || (xpc10nz==9'd451/*451:US*/) || (xpc10nz==9'd457/*457:US*/) || (xpc10nz==9'd478/*478:US*/)) && 
              !xpc10_stall;

               Z64SSCCSCALbx54ARB0RRh10shot0 <= ((TSPcr2_16_V_1<32'd77) && (xpc10nz==9'd461/*461:US*/) || (xpc10nz==9'd424/*424:US*/) || 
              (xpc10nz==9'd413/*413:US*/) || (xpc10nz==9'd444/*444:US*/)) && !xpc10_stall;

               iuMULTIPLIER14RRh12shot0 <= ((TSPcr2_16_V_1<32'd77) && (xpc10nz==9'd459/*459:US*/) || (xpc10nz==9'd436/*436:US*/) || (xpc10nz
              ==9'd426/*426:US*/) || (xpc10nz==9'd416/*416:US*/) || (xpc10nz==9'd403/*403:US*/) || (xpc10nz==9'd411/*411:US*/) || (xpc10nz
              ==9'd422/*422:US*/) || (xpc10nz==9'd430/*430:US*/) || (xpc10nz==9'd442/*442:US*/)) && !xpc10_stall;

               Z64SSCCSCALbx58ARD0RRh10shot0 <= ((xpc10nz==9'd438/*438:US*/) || (xpc10nz==9'd428/*428:US*/)) && !xpc10_stall;
               Z64SSCCSCALbx52ARA0RRh10shot0 <= ((xpc10nz==9'd438/*438:US*/) || (xpc10nz==9'd432/*432:US*/)) && !xpc10_stall;
               iuMULTIPLIER12RRh10shot0 <= ((xpc10nz==9'd436/*436:US*/) || (xpc10nz==9'd426/*426:US*/) || (xpc10nz==9'd402/*402:US*/) || 
              (xpc10nz==9'd411/*411:US*/) || (xpc10nz==9'd430/*430:US*/)) && !xpc10_stall;

               Z64SSCCSCALbx56ARC0RRh10shot0 <= ((xpc10nz==9'd432/*432:US*/) || (xpc10nz==9'd428/*428:US*/)) && !xpc10_stall;
               SINTCCSCALbx16ARA0RRh10shot0 <= (xpc10nz==9'd418/*418:US*/) && !xpc10_stall;
               Z16SSCCSCALbx10ARA0RRh10shot0 <= (xpc10nz==9'd409/*409:US*/) && !xpc10_stall;
               iuMULTIPLIER14RRh10shot0 <= (xpc10nz==9'd402/*402:US*/) && !xpc10_stall;
               iuMULTIPLIER10RRh10shot0 <= (xpc10nz==9'd402/*402:US*/) && !xpc10_stall;
              if ((xpc10nz==1'd1/*1:US*/))  xpc10nz <= 2'd2/*2:xpc10nz*/;
                  if ((xpc10nz==2'd2/*2:US*/))  xpc10nz <= 2'd3/*3:xpc10nz*/;
                  if ((xpc10nz==2'd3/*3:US*/))  xpc10nz <= 3'd4/*4:xpc10nz*/;
                  if ((xpc10nz==3'd4/*4:US*/))  xpc10nz <= 3'd5/*5:xpc10nz*/;
                  if ((xpc10nz==3'd5/*5:US*/))  xpc10nz <= 3'd6/*6:xpc10nz*/;
                  if ((xpc10nz==3'd6/*6:US*/))  xpc10nz <= 3'd7/*7:xpc10nz*/;
                  if ((xpc10nz==3'd7/*7:US*/))  xpc10nz <= 4'd8/*8:xpc10nz*/;
                  if ((xpc10nz==4'd8/*8:US*/))  xpc10nz <= 4'd9/*9:xpc10nz*/;
                  if ((xpc10nz==4'd9/*9:US*/))  xpc10nz <= 4'd10/*10:xpc10nz*/;
                  if ((xpc10nz==4'd10/*10:US*/))  xpc10nz <= 4'd11/*11:xpc10nz*/;
                  if ((xpc10nz==4'd11/*11:US*/))  xpc10nz <= 4'd12/*12:xpc10nz*/;
                  if ((xpc10nz==4'd12/*12:US*/))  xpc10nz <= 4'd13/*13:xpc10nz*/;
                  if ((xpc10nz==4'd13/*13:US*/))  xpc10nz <= 4'd14/*14:xpc10nz*/;
                  if ((xpc10nz==4'd14/*14:US*/))  xpc10nz <= 4'd15/*15:xpc10nz*/;
                  if ((xpc10nz==4'd15/*15:US*/))  xpc10nz <= 5'd16/*16:xpc10nz*/;
                  if ((xpc10nz==5'd16/*16:US*/))  xpc10nz <= 5'd17/*17:xpc10nz*/;
                  if ((xpc10nz==5'd17/*17:US*/))  xpc10nz <= 5'd18/*18:xpc10nz*/;
                  if ((xpc10nz==5'd18/*18:US*/))  xpc10nz <= 5'd19/*19:xpc10nz*/;
                  if ((xpc10nz==5'd19/*19:US*/))  xpc10nz <= 5'd20/*20:xpc10nz*/;
                  if ((xpc10nz==5'd20/*20:US*/))  xpc10nz <= 5'd21/*21:xpc10nz*/;
                  if ((xpc10nz==5'd21/*21:US*/))  xpc10nz <= 5'd22/*22:xpc10nz*/;
                  if ((xpc10nz==5'd22/*22:US*/))  xpc10nz <= 5'd23/*23:xpc10nz*/;
                  if ((xpc10nz==5'd23/*23:US*/))  xpc10nz <= 5'd24/*24:xpc10nz*/;
                  if ((xpc10nz==5'd24/*24:US*/))  xpc10nz <= 5'd25/*25:xpc10nz*/;
                  if ((xpc10nz==5'd25/*25:US*/))  xpc10nz <= 5'd26/*26:xpc10nz*/;
                  if ((xpc10nz==5'd26/*26:US*/))  xpc10nz <= 5'd27/*27:xpc10nz*/;
                  if ((xpc10nz==5'd27/*27:US*/))  xpc10nz <= 5'd28/*28:xpc10nz*/;
                  if ((xpc10nz==5'd28/*28:US*/))  xpc10nz <= 5'd29/*29:xpc10nz*/;
                  if ((xpc10nz==5'd29/*29:US*/))  xpc10nz <= 5'd30/*30:xpc10nz*/;
                  if ((xpc10nz==5'd30/*30:US*/))  xpc10nz <= 5'd31/*31:xpc10nz*/;
                  if ((xpc10nz==5'd31/*31:US*/))  xpc10nz <= 6'd32/*32:xpc10nz*/;
                  if ((xpc10nz==6'd32/*32:US*/))  xpc10nz <= 6'd33/*33:xpc10nz*/;
                  if ((xpc10nz==6'd33/*33:US*/))  xpc10nz <= 6'd34/*34:xpc10nz*/;
                  if ((xpc10nz==6'd34/*34:US*/))  xpc10nz <= 6'd35/*35:xpc10nz*/;
                  if ((xpc10nz==6'd35/*35:US*/))  xpc10nz <= 6'd36/*36:xpc10nz*/;
                  if ((xpc10nz==6'd36/*36:US*/))  xpc10nz <= 6'd37/*37:xpc10nz*/;
                  if ((xpc10nz==6'd37/*37:US*/))  xpc10nz <= 6'd38/*38:xpc10nz*/;
                  if ((xpc10nz==6'd38/*38:US*/))  xpc10nz <= 6'd39/*39:xpc10nz*/;
                  if ((xpc10nz==6'd39/*39:US*/))  xpc10nz <= 6'd40/*40:xpc10nz*/;
                  if ((xpc10nz==6'd40/*40:US*/))  xpc10nz <= 6'd41/*41:xpc10nz*/;
                  if ((xpc10nz==6'd41/*41:US*/))  xpc10nz <= 6'd42/*42:xpc10nz*/;
                  if ((xpc10nz==6'd42/*42:US*/))  xpc10nz <= 6'd43/*43:xpc10nz*/;
                  if ((xpc10nz==6'd43/*43:US*/))  xpc10nz <= 6'd44/*44:xpc10nz*/;
                  if ((xpc10nz==6'd44/*44:US*/))  xpc10nz <= 6'd45/*45:xpc10nz*/;
                  if ((xpc10nz==6'd45/*45:US*/))  xpc10nz <= 6'd46/*46:xpc10nz*/;
                  if ((xpc10nz==6'd46/*46:US*/))  xpc10nz <= 6'd47/*47:xpc10nz*/;
                  if ((xpc10nz==6'd47/*47:US*/))  xpc10nz <= 6'd48/*48:xpc10nz*/;
                  if ((xpc10nz==6'd48/*48:US*/))  xpc10nz <= 6'd49/*49:xpc10nz*/;
                  if ((xpc10nz==6'd49/*49:US*/))  xpc10nz <= 6'd50/*50:xpc10nz*/;
                  if ((xpc10nz==6'd50/*50:US*/))  xpc10nz <= 6'd51/*51:xpc10nz*/;
                  if ((xpc10nz==6'd51/*51:US*/))  xpc10nz <= 6'd52/*52:xpc10nz*/;
                  if ((xpc10nz==6'd52/*52:US*/))  xpc10nz <= 6'd53/*53:xpc10nz*/;
                  if ((xpc10nz==6'd53/*53:US*/))  xpc10nz <= 6'd54/*54:xpc10nz*/;
                  if ((xpc10nz==6'd54/*54:US*/))  xpc10nz <= 6'd55/*55:xpc10nz*/;
                  if ((xpc10nz==6'd55/*55:US*/))  xpc10nz <= 6'd56/*56:xpc10nz*/;
                  if ((xpc10nz==6'd56/*56:US*/))  xpc10nz <= 6'd57/*57:xpc10nz*/;
                  if ((xpc10nz==6'd57/*57:US*/))  xpc10nz <= 6'd58/*58:xpc10nz*/;
                  if ((xpc10nz==6'd58/*58:US*/))  xpc10nz <= 6'd59/*59:xpc10nz*/;
                  if ((xpc10nz==6'd59/*59:US*/))  xpc10nz <= 6'd60/*60:xpc10nz*/;
                  if ((xpc10nz==6'd60/*60:US*/))  xpc10nz <= 6'd61/*61:xpc10nz*/;
                  if ((xpc10nz==6'd61/*61:US*/))  xpc10nz <= 6'd62/*62:xpc10nz*/;
                  if ((xpc10nz==6'd62/*62:US*/))  xpc10nz <= 6'd63/*63:xpc10nz*/;
                  if ((xpc10nz==6'd63/*63:US*/))  xpc10nz <= 7'd64/*64:xpc10nz*/;
                  if ((xpc10nz==7'd64/*64:US*/))  xpc10nz <= 7'd65/*65:xpc10nz*/;
                  if ((xpc10nz==7'd65/*65:US*/))  xpc10nz <= 7'd66/*66:xpc10nz*/;
                  if ((xpc10nz==7'd66/*66:US*/))  xpc10nz <= 7'd67/*67:xpc10nz*/;
                  if ((xpc10nz==7'd67/*67:US*/))  xpc10nz <= 7'd68/*68:xpc10nz*/;
                  if ((xpc10nz==7'd68/*68:US*/))  xpc10nz <= 7'd69/*69:xpc10nz*/;
                  if ((xpc10nz==7'd69/*69:US*/))  xpc10nz <= 7'd70/*70:xpc10nz*/;
                  if ((xpc10nz==7'd70/*70:US*/))  xpc10nz <= 7'd71/*71:xpc10nz*/;
                  if ((xpc10nz==7'd71/*71:US*/))  xpc10nz <= 7'd72/*72:xpc10nz*/;
                  if ((xpc10nz==7'd72/*72:US*/))  xpc10nz <= 7'd73/*73:xpc10nz*/;
                  if ((xpc10nz==7'd73/*73:US*/))  xpc10nz <= 7'd74/*74:xpc10nz*/;
                  if ((xpc10nz==7'd74/*74:US*/))  xpc10nz <= 7'd75/*75:xpc10nz*/;
                  if ((xpc10nz==7'd75/*75:US*/))  xpc10nz <= 7'd76/*76:xpc10nz*/;
                  if ((xpc10nz==7'd76/*76:US*/))  xpc10nz <= 7'd77/*77:xpc10nz*/;
                  if ((xpc10nz==7'd77/*77:US*/))  xpc10nz <= 7'd78/*78:xpc10nz*/;
                  if ((xpc10nz==7'd78/*78:US*/))  xpc10nz <= 7'd79/*79:xpc10nz*/;
                  if ((xpc10nz==7'd79/*79:US*/))  xpc10nz <= 7'd80/*80:xpc10nz*/;
                  if ((xpc10nz==7'd80/*80:US*/))  xpc10nz <= 7'd81/*81:xpc10nz*/;
                  if ((xpc10nz==7'd81/*81:US*/))  xpc10nz <= 7'd82/*82:xpc10nz*/;
                  if ((xpc10nz==7'd82/*82:US*/))  xpc10nz <= 7'd83/*83:xpc10nz*/;
                  if ((xpc10nz==7'd83/*83:US*/))  xpc10nz <= 7'd84/*84:xpc10nz*/;
                  if ((xpc10nz==7'd84/*84:US*/))  xpc10nz <= 7'd85/*85:xpc10nz*/;
                  if ((xpc10nz==7'd85/*85:US*/))  xpc10nz <= 7'd86/*86:xpc10nz*/;
                  if ((xpc10nz==7'd86/*86:US*/))  xpc10nz <= 7'd87/*87:xpc10nz*/;
                  if ((xpc10nz==7'd87/*87:US*/))  xpc10nz <= 7'd88/*88:xpc10nz*/;
                  if ((xpc10nz==7'd88/*88:US*/))  xpc10nz <= 7'd89/*89:xpc10nz*/;
                  if ((xpc10nz==7'd89/*89:US*/))  xpc10nz <= 7'd90/*90:xpc10nz*/;
                  if ((xpc10nz==7'd90/*90:US*/))  xpc10nz <= 7'd91/*91:xpc10nz*/;
                  if ((xpc10nz==7'd91/*91:US*/))  xpc10nz <= 7'd92/*92:xpc10nz*/;
                  if ((xpc10nz==7'd92/*92:US*/))  xpc10nz <= 7'd93/*93:xpc10nz*/;
                  if ((xpc10nz==7'd93/*93:US*/))  xpc10nz <= 7'd94/*94:xpc10nz*/;
                  if ((xpc10nz==7'd94/*94:US*/))  xpc10nz <= 7'd95/*95:xpc10nz*/;
                  if ((xpc10nz==7'd95/*95:US*/))  xpc10nz <= 7'd96/*96:xpc10nz*/;
                  if ((xpc10nz==7'd96/*96:US*/))  xpc10nz <= 7'd97/*97:xpc10nz*/;
                  if ((xpc10nz==7'd97/*97:US*/))  xpc10nz <= 7'd98/*98:xpc10nz*/;
                  if ((xpc10nz==7'd98/*98:US*/))  xpc10nz <= 7'd99/*99:xpc10nz*/;
                  if ((xpc10nz==7'd99/*99:US*/))  xpc10nz <= 7'd100/*100:xpc10nz*/;
                  if ((xpc10nz==7'd100/*100:US*/))  xpc10nz <= 7'd101/*101:xpc10nz*/;
                  if ((xpc10nz==7'd101/*101:US*/))  xpc10nz <= 7'd102/*102:xpc10nz*/;
                  if ((xpc10nz==7'd102/*102:US*/))  xpc10nz <= 7'd103/*103:xpc10nz*/;
                  if ((xpc10nz==7'd103/*103:US*/))  xpc10nz <= 7'd104/*104:xpc10nz*/;
                  if ((xpc10nz==7'd104/*104:US*/))  xpc10nz <= 7'd105/*105:xpc10nz*/;
                  if ((xpc10nz==7'd105/*105:US*/))  xpc10nz <= 7'd106/*106:xpc10nz*/;
                  if ((xpc10nz==7'd106/*106:US*/))  xpc10nz <= 7'd107/*107:xpc10nz*/;
                  if ((xpc10nz==7'd107/*107:US*/))  xpc10nz <= 7'd108/*108:xpc10nz*/;
                  if ((xpc10nz==7'd108/*108:US*/))  xpc10nz <= 7'd109/*109:xpc10nz*/;
                  if ((xpc10nz==7'd109/*109:US*/))  xpc10nz <= 7'd110/*110:xpc10nz*/;
                  if ((xpc10nz==7'd110/*110:US*/))  xpc10nz <= 7'd111/*111:xpc10nz*/;
                  if ((xpc10nz==7'd111/*111:US*/))  xpc10nz <= 7'd112/*112:xpc10nz*/;
                  if ((xpc10nz==7'd112/*112:US*/))  xpc10nz <= 7'd113/*113:xpc10nz*/;
                  if ((xpc10nz==7'd113/*113:US*/))  xpc10nz <= 7'd114/*114:xpc10nz*/;
                  if ((xpc10nz==7'd114/*114:US*/))  xpc10nz <= 7'd115/*115:xpc10nz*/;
                  if ((xpc10nz==7'd115/*115:US*/))  xpc10nz <= 7'd116/*116:xpc10nz*/;
                  if ((xpc10nz==7'd116/*116:US*/))  xpc10nz <= 7'd117/*117:xpc10nz*/;
                  if ((xpc10nz==7'd117/*117:US*/))  xpc10nz <= 7'd118/*118:xpc10nz*/;
                  if ((xpc10nz==7'd118/*118:US*/))  xpc10nz <= 7'd119/*119:xpc10nz*/;
                  if ((xpc10nz==7'd119/*119:US*/))  xpc10nz <= 7'd120/*120:xpc10nz*/;
                  if ((xpc10nz==7'd120/*120:US*/))  xpc10nz <= 7'd121/*121:xpc10nz*/;
                  if ((xpc10nz==7'd121/*121:US*/))  xpc10nz <= 7'd122/*122:xpc10nz*/;
                  if ((xpc10nz==7'd122/*122:US*/))  xpc10nz <= 7'd123/*123:xpc10nz*/;
                  if ((xpc10nz==7'd123/*123:US*/))  xpc10nz <= 7'd124/*124:xpc10nz*/;
                  if ((xpc10nz==7'd124/*124:US*/))  xpc10nz <= 7'd125/*125:xpc10nz*/;
                  if ((xpc10nz==7'd125/*125:US*/))  xpc10nz <= 7'd126/*126:xpc10nz*/;
                  if ((xpc10nz==7'd126/*126:US*/))  xpc10nz <= 7'd127/*127:xpc10nz*/;
                  if ((xpc10nz==7'd127/*127:US*/))  xpc10nz <= 8'd128/*128:xpc10nz*/;
                  if ((xpc10nz==8'd128/*128:US*/))  xpc10nz <= 8'd129/*129:xpc10nz*/;
                  if ((xpc10nz==8'd129/*129:US*/))  xpc10nz <= 8'd130/*130:xpc10nz*/;
                  if ((xpc10nz==8'd130/*130:US*/))  xpc10nz <= 8'd131/*131:xpc10nz*/;
                  if ((xpc10nz==8'd131/*131:US*/))  xpc10nz <= 8'd132/*132:xpc10nz*/;
                  if ((xpc10nz==8'd132/*132:US*/))  xpc10nz <= 8'd133/*133:xpc10nz*/;
                  if ((xpc10nz==8'd133/*133:US*/))  xpc10nz <= 8'd134/*134:xpc10nz*/;
                  if ((xpc10nz==8'd134/*134:US*/))  xpc10nz <= 8'd135/*135:xpc10nz*/;
                  if ((xpc10nz==8'd135/*135:US*/))  xpc10nz <= 8'd136/*136:xpc10nz*/;
                  if ((xpc10nz==8'd136/*136:US*/))  xpc10nz <= 8'd137/*137:xpc10nz*/;
                  if ((xpc10nz==8'd137/*137:US*/))  xpc10nz <= 8'd138/*138:xpc10nz*/;
                  if ((xpc10nz==8'd138/*138:US*/))  xpc10nz <= 8'd139/*139:xpc10nz*/;
                  if ((xpc10nz==8'd139/*139:US*/))  xpc10nz <= 8'd140/*140:xpc10nz*/;
                  if ((xpc10nz==8'd140/*140:US*/))  xpc10nz <= 8'd141/*141:xpc10nz*/;
                  if ((xpc10nz==8'd141/*141:US*/))  xpc10nz <= 8'd142/*142:xpc10nz*/;
                  if ((xpc10nz==8'd142/*142:US*/))  xpc10nz <= 8'd143/*143:xpc10nz*/;
                  if ((xpc10nz==8'd143/*143:US*/))  xpc10nz <= 8'd144/*144:xpc10nz*/;
                  if ((xpc10nz==8'd144/*144:US*/))  xpc10nz <= 8'd145/*145:xpc10nz*/;
                  if ((xpc10nz==8'd145/*145:US*/))  xpc10nz <= 8'd146/*146:xpc10nz*/;
                  if ((xpc10nz==8'd146/*146:US*/))  xpc10nz <= 8'd147/*147:xpc10nz*/;
                  if ((xpc10nz==8'd147/*147:US*/))  xpc10nz <= 8'd148/*148:xpc10nz*/;
                  if ((xpc10nz==8'd148/*148:US*/))  xpc10nz <= 8'd149/*149:xpc10nz*/;
                  if ((xpc10nz==8'd149/*149:US*/))  xpc10nz <= 8'd150/*150:xpc10nz*/;
                  if ((xpc10nz==8'd150/*150:US*/))  xpc10nz <= 8'd151/*151:xpc10nz*/;
                  if ((xpc10nz==8'd151/*151:US*/))  xpc10nz <= 8'd152/*152:xpc10nz*/;
                  if ((xpc10nz==8'd152/*152:US*/))  xpc10nz <= 8'd153/*153:xpc10nz*/;
                  if ((xpc10nz==8'd153/*153:US*/))  xpc10nz <= 8'd154/*154:xpc10nz*/;
                  if ((xpc10nz==8'd154/*154:US*/))  xpc10nz <= 8'd155/*155:xpc10nz*/;
                  if ((xpc10nz==8'd155/*155:US*/))  xpc10nz <= 8'd156/*156:xpc10nz*/;
                  if ((xpc10nz==8'd156/*156:US*/))  xpc10nz <= 8'd157/*157:xpc10nz*/;
                  if ((xpc10nz==8'd157/*157:US*/))  xpc10nz <= 8'd158/*158:xpc10nz*/;
                  if ((xpc10nz==8'd158/*158:US*/))  xpc10nz <= 8'd159/*159:xpc10nz*/;
                  if ((xpc10nz==8'd159/*159:US*/))  xpc10nz <= 8'd160/*160:xpc10nz*/;
                  if ((xpc10nz==8'd160/*160:US*/))  xpc10nz <= 8'd161/*161:xpc10nz*/;
                  if ((xpc10nz==8'd161/*161:US*/))  xpc10nz <= 8'd162/*162:xpc10nz*/;
                  if ((xpc10nz==8'd162/*162:US*/))  xpc10nz <= 8'd163/*163:xpc10nz*/;
                  if ((xpc10nz==8'd163/*163:US*/))  xpc10nz <= 8'd164/*164:xpc10nz*/;
                  if ((xpc10nz==8'd164/*164:US*/))  xpc10nz <= 8'd165/*165:xpc10nz*/;
                  if ((xpc10nz==8'd165/*165:US*/))  xpc10nz <= 8'd166/*166:xpc10nz*/;
                  if ((xpc10nz==8'd166/*166:US*/))  xpc10nz <= 8'd167/*167:xpc10nz*/;
                  if ((xpc10nz==8'd167/*167:US*/))  xpc10nz <= 8'd168/*168:xpc10nz*/;
                  if ((xpc10nz==8'd168/*168:US*/))  xpc10nz <= 8'd169/*169:xpc10nz*/;
                  if ((xpc10nz==8'd169/*169:US*/))  xpc10nz <= 8'd170/*170:xpc10nz*/;
                  if ((xpc10nz==8'd170/*170:US*/))  xpc10nz <= 8'd171/*171:xpc10nz*/;
                  if ((xpc10nz==8'd171/*171:US*/))  xpc10nz <= 8'd172/*172:xpc10nz*/;
                  if ((xpc10nz==8'd172/*172:US*/))  xpc10nz <= 8'd173/*173:xpc10nz*/;
                  if ((xpc10nz==8'd173/*173:US*/))  xpc10nz <= 8'd174/*174:xpc10nz*/;
                  if ((xpc10nz==8'd174/*174:US*/))  xpc10nz <= 8'd175/*175:xpc10nz*/;
                  if ((xpc10nz==8'd175/*175:US*/))  xpc10nz <= 8'd176/*176:xpc10nz*/;
                  if ((xpc10nz==8'd176/*176:US*/))  xpc10nz <= 8'd177/*177:xpc10nz*/;
                  if ((xpc10nz==8'd177/*177:US*/))  xpc10nz <= 8'd178/*178:xpc10nz*/;
                  if ((xpc10nz==8'd178/*178:US*/))  xpc10nz <= 8'd179/*179:xpc10nz*/;
                  if ((xpc10nz==8'd179/*179:US*/))  xpc10nz <= 8'd180/*180:xpc10nz*/;
                  if ((xpc10nz==8'd180/*180:US*/))  xpc10nz <= 8'd181/*181:xpc10nz*/;
                  if ((xpc10nz==8'd181/*181:US*/))  xpc10nz <= 8'd182/*182:xpc10nz*/;
                  if ((xpc10nz==8'd182/*182:US*/))  xpc10nz <= 8'd183/*183:xpc10nz*/;
                  if ((xpc10nz==8'd183/*183:US*/))  xpc10nz <= 8'd184/*184:xpc10nz*/;
                  if ((xpc10nz==8'd184/*184:US*/))  xpc10nz <= 8'd185/*185:xpc10nz*/;
                  if ((xpc10nz==8'd185/*185:US*/))  xpc10nz <= 8'd186/*186:xpc10nz*/;
                  if ((xpc10nz==8'd186/*186:US*/))  xpc10nz <= 8'd187/*187:xpc10nz*/;
                  if ((xpc10nz==8'd187/*187:US*/))  xpc10nz <= 8'd188/*188:xpc10nz*/;
                  if ((xpc10nz==8'd188/*188:US*/))  xpc10nz <= 8'd189/*189:xpc10nz*/;
                  if ((xpc10nz==8'd189/*189:US*/))  xpc10nz <= 8'd190/*190:xpc10nz*/;
                  if ((xpc10nz==8'd190/*190:US*/))  xpc10nz <= 8'd191/*191:xpc10nz*/;
                  if ((xpc10nz==8'd191/*191:US*/))  xpc10nz <= 8'd192/*192:xpc10nz*/;
                  if ((xpc10nz==8'd192/*192:US*/))  xpc10nz <= 8'd193/*193:xpc10nz*/;
                  if ((xpc10nz==8'd193/*193:US*/))  xpc10nz <= 8'd194/*194:xpc10nz*/;
                  if ((xpc10nz==8'd194/*194:US*/))  xpc10nz <= 8'd195/*195:xpc10nz*/;
                  if ((xpc10nz==8'd195/*195:US*/))  xpc10nz <= 8'd196/*196:xpc10nz*/;
                  if ((xpc10nz==8'd196/*196:US*/))  xpc10nz <= 8'd197/*197:xpc10nz*/;
                  if ((xpc10nz==8'd197/*197:US*/))  xpc10nz <= 8'd198/*198:xpc10nz*/;
                  if ((xpc10nz==8'd198/*198:US*/))  xpc10nz <= 8'd199/*199:xpc10nz*/;
                  if ((xpc10nz==8'd199/*199:US*/))  xpc10nz <= 8'd200/*200:xpc10nz*/;
                  if ((xpc10nz==8'd200/*200:US*/))  xpc10nz <= 8'd201/*201:xpc10nz*/;
                  if ((xpc10nz==8'd201/*201:US*/))  xpc10nz <= 8'd202/*202:xpc10nz*/;
                  if ((xpc10nz==8'd202/*202:US*/))  xpc10nz <= 8'd203/*203:xpc10nz*/;
                  if ((xpc10nz==8'd203/*203:US*/))  xpc10nz <= 8'd204/*204:xpc10nz*/;
                  if ((xpc10nz==8'd204/*204:US*/))  xpc10nz <= 8'd205/*205:xpc10nz*/;
                  if ((xpc10nz==8'd205/*205:US*/))  xpc10nz <= 8'd206/*206:xpc10nz*/;
                  if ((xpc10nz==8'd206/*206:US*/))  xpc10nz <= 8'd207/*207:xpc10nz*/;
                  if ((xpc10nz==8'd207/*207:US*/))  xpc10nz <= 8'd208/*208:xpc10nz*/;
                  if ((xpc10nz==8'd208/*208:US*/))  xpc10nz <= 8'd209/*209:xpc10nz*/;
                  if ((xpc10nz==8'd209/*209:US*/))  xpc10nz <= 8'd210/*210:xpc10nz*/;
                  if ((xpc10nz==8'd210/*210:US*/))  xpc10nz <= 8'd211/*211:xpc10nz*/;
                  if ((xpc10nz==8'd211/*211:US*/))  xpc10nz <= 8'd212/*212:xpc10nz*/;
                  if ((xpc10nz==8'd212/*212:US*/))  xpc10nz <= 8'd213/*213:xpc10nz*/;
                  if ((xpc10nz==8'd213/*213:US*/))  xpc10nz <= 8'd214/*214:xpc10nz*/;
                  if ((xpc10nz==8'd214/*214:US*/))  xpc10nz <= 8'd215/*215:xpc10nz*/;
                  if ((xpc10nz==8'd215/*215:US*/))  xpc10nz <= 8'd216/*216:xpc10nz*/;
                  if ((xpc10nz==8'd216/*216:US*/))  xpc10nz <= 8'd217/*217:xpc10nz*/;
                  if ((xpc10nz==8'd217/*217:US*/))  xpc10nz <= 8'd218/*218:xpc10nz*/;
                  if ((xpc10nz==8'd218/*218:US*/))  xpc10nz <= 8'd219/*219:xpc10nz*/;
                  if ((xpc10nz==8'd219/*219:US*/))  xpc10nz <= 8'd220/*220:xpc10nz*/;
                  if ((xpc10nz==8'd220/*220:US*/))  xpc10nz <= 8'd221/*221:xpc10nz*/;
                  if ((xpc10nz==8'd221/*221:US*/))  xpc10nz <= 8'd222/*222:xpc10nz*/;
                  if ((xpc10nz==8'd222/*222:US*/))  xpc10nz <= 8'd223/*223:xpc10nz*/;
                  if ((xpc10nz==8'd223/*223:US*/))  xpc10nz <= 8'd224/*224:xpc10nz*/;
                  if ((xpc10nz==8'd224/*224:US*/))  xpc10nz <= 8'd225/*225:xpc10nz*/;
                  if ((xpc10nz==8'd225/*225:US*/))  xpc10nz <= 8'd226/*226:xpc10nz*/;
                  if ((xpc10nz==8'd226/*226:US*/))  xpc10nz <= 8'd227/*227:xpc10nz*/;
                  if ((xpc10nz==8'd227/*227:US*/))  xpc10nz <= 8'd228/*228:xpc10nz*/;
                  if ((xpc10nz==8'd228/*228:US*/))  xpc10nz <= 8'd229/*229:xpc10nz*/;
                  if ((xpc10nz==8'd229/*229:US*/))  xpc10nz <= 8'd230/*230:xpc10nz*/;
                  if ((xpc10nz==8'd230/*230:US*/))  xpc10nz <= 8'd231/*231:xpc10nz*/;
                  if ((xpc10nz==8'd231/*231:US*/))  xpc10nz <= 8'd232/*232:xpc10nz*/;
                  if ((xpc10nz==8'd232/*232:US*/))  xpc10nz <= 8'd233/*233:xpc10nz*/;
                  if ((xpc10nz==8'd233/*233:US*/))  xpc10nz <= 8'd234/*234:xpc10nz*/;
                  if ((xpc10nz==8'd234/*234:US*/))  xpc10nz <= 8'd235/*235:xpc10nz*/;
                  if ((xpc10nz==8'd235/*235:US*/))  xpc10nz <= 8'd236/*236:xpc10nz*/;
                  if ((xpc10nz==8'd236/*236:US*/))  xpc10nz <= 8'd237/*237:xpc10nz*/;
                  if ((xpc10nz==8'd237/*237:US*/))  xpc10nz <= 8'd238/*238:xpc10nz*/;
                  if ((xpc10nz==8'd238/*238:US*/))  xpc10nz <= 8'd239/*239:xpc10nz*/;
                  if ((xpc10nz==8'd239/*239:US*/))  xpc10nz <= 8'd240/*240:xpc10nz*/;
                  if ((xpc10nz==8'd240/*240:US*/))  xpc10nz <= 8'd241/*241:xpc10nz*/;
                  if ((xpc10nz==8'd241/*241:US*/))  xpc10nz <= 8'd242/*242:xpc10nz*/;
                  if ((xpc10nz==8'd242/*242:US*/))  xpc10nz <= 8'd243/*243:xpc10nz*/;
                  if ((xpc10nz==8'd243/*243:US*/))  xpc10nz <= 8'd244/*244:xpc10nz*/;
                  if ((xpc10nz==8'd244/*244:US*/))  xpc10nz <= 8'd245/*245:xpc10nz*/;
                  if ((xpc10nz==8'd245/*245:US*/))  xpc10nz <= 8'd246/*246:xpc10nz*/;
                  if ((xpc10nz==8'd246/*246:US*/))  xpc10nz <= 8'd247/*247:xpc10nz*/;
                  if ((xpc10nz==8'd247/*247:US*/))  xpc10nz <= 8'd248/*248:xpc10nz*/;
                  if ((xpc10nz==8'd248/*248:US*/))  xpc10nz <= 8'd249/*249:xpc10nz*/;
                  if ((xpc10nz==8'd249/*249:US*/))  xpc10nz <= 8'd250/*250:xpc10nz*/;
                  if ((xpc10nz==8'd250/*250:US*/))  xpc10nz <= 8'd251/*251:xpc10nz*/;
                  if ((xpc10nz==8'd251/*251:US*/))  xpc10nz <= 8'd252/*252:xpc10nz*/;
                  if ((xpc10nz==8'd252/*252:US*/))  xpc10nz <= 8'd253/*253:xpc10nz*/;
                  if ((xpc10nz==8'd253/*253:US*/))  xpc10nz <= 8'd254/*254:xpc10nz*/;
                  if ((xpc10nz==8'd254/*254:US*/))  xpc10nz <= 8'd255/*255:xpc10nz*/;
                  if ((xpc10nz==8'd255/*255:US*/))  xpc10nz <= 9'd256/*256:xpc10nz*/;
                  if ((xpc10nz==9'd256/*256:US*/))  xpc10nz <= 9'd257/*257:xpc10nz*/;
                  if ((xpc10nz==9'd257/*257:US*/))  xpc10nz <= 9'd258/*258:xpc10nz*/;
                  if ((xpc10nz==9'd258/*258:US*/))  xpc10nz <= 9'd259/*259:xpc10nz*/;
                  if ((xpc10nz==9'd259/*259:US*/))  xpc10nz <= 9'd260/*260:xpc10nz*/;
                  if ((xpc10nz==9'd260/*260:US*/))  xpc10nz <= 9'd261/*261:xpc10nz*/;
                  if ((xpc10nz==9'd261/*261:US*/))  xpc10nz <= 9'd262/*262:xpc10nz*/;
                  if ((xpc10nz==9'd262/*262:US*/))  xpc10nz <= 9'd263/*263:xpc10nz*/;
                  if ((xpc10nz==9'd263/*263:US*/))  xpc10nz <= 9'd264/*264:xpc10nz*/;
                  if ((xpc10nz==9'd264/*264:US*/))  xpc10nz <= 9'd265/*265:xpc10nz*/;
                  if ((xpc10nz==9'd265/*265:US*/))  xpc10nz <= 9'd266/*266:xpc10nz*/;
                  if ((xpc10nz==9'd266/*266:US*/))  xpc10nz <= 9'd267/*267:xpc10nz*/;
                  if ((xpc10nz==9'd267/*267:US*/))  xpc10nz <= 9'd268/*268:xpc10nz*/;
                  if ((xpc10nz==9'd268/*268:US*/))  xpc10nz <= 9'd269/*269:xpc10nz*/;
                  if ((xpc10nz==9'd269/*269:US*/))  xpc10nz <= 9'd270/*270:xpc10nz*/;
                  if ((xpc10nz==9'd270/*270:US*/))  xpc10nz <= 9'd271/*271:xpc10nz*/;
                  if ((xpc10nz==9'd271/*271:US*/))  xpc10nz <= 9'd272/*272:xpc10nz*/;
                  if ((xpc10nz==9'd272/*272:US*/))  xpc10nz <= 9'd273/*273:xpc10nz*/;
                  if ((xpc10nz==9'd273/*273:US*/))  xpc10nz <= 9'd274/*274:xpc10nz*/;
                  if ((xpc10nz==9'd274/*274:US*/))  xpc10nz <= 9'd275/*275:xpc10nz*/;
                  if ((xpc10nz==9'd275/*275:US*/))  xpc10nz <= 9'd276/*276:xpc10nz*/;
                  if ((xpc10nz==9'd276/*276:US*/))  xpc10nz <= 9'd277/*277:xpc10nz*/;
                  if ((xpc10nz==9'd277/*277:US*/))  xpc10nz <= 9'd278/*278:xpc10nz*/;
                  if ((xpc10nz==9'd278/*278:US*/))  xpc10nz <= 9'd279/*279:xpc10nz*/;
                  if ((xpc10nz==9'd279/*279:US*/))  xpc10nz <= 9'd280/*280:xpc10nz*/;
                  if ((xpc10nz==9'd280/*280:US*/))  xpc10nz <= 9'd281/*281:xpc10nz*/;
                  if ((xpc10nz==9'd281/*281:US*/))  xpc10nz <= 9'd282/*282:xpc10nz*/;
                  if ((xpc10nz==9'd282/*282:US*/))  xpc10nz <= 9'd283/*283:xpc10nz*/;
                  if ((xpc10nz==9'd283/*283:US*/))  xpc10nz <= 9'd284/*284:xpc10nz*/;
                  if ((xpc10nz==9'd284/*284:US*/))  xpc10nz <= 9'd285/*285:xpc10nz*/;
                  if ((xpc10nz==9'd285/*285:US*/))  xpc10nz <= 9'd286/*286:xpc10nz*/;
                  if ((xpc10nz==9'd286/*286:US*/))  xpc10nz <= 9'd287/*287:xpc10nz*/;
                  if ((xpc10nz==9'd287/*287:US*/))  xpc10nz <= 9'd288/*288:xpc10nz*/;
                  if ((xpc10nz==9'd288/*288:US*/))  xpc10nz <= 9'd289/*289:xpc10nz*/;
                  if ((xpc10nz==9'd289/*289:US*/))  xpc10nz <= 9'd290/*290:xpc10nz*/;
                  if ((xpc10nz==9'd290/*290:US*/))  xpc10nz <= 9'd291/*291:xpc10nz*/;
                  if ((xpc10nz==9'd291/*291:US*/))  xpc10nz <= 9'd292/*292:xpc10nz*/;
                  if ((xpc10nz==9'd292/*292:US*/))  xpc10nz <= 9'd293/*293:xpc10nz*/;
                  if ((xpc10nz==9'd293/*293:US*/))  xpc10nz <= 9'd294/*294:xpc10nz*/;
                  if ((xpc10nz==9'd294/*294:US*/))  xpc10nz <= 9'd295/*295:xpc10nz*/;
                  if ((xpc10nz==9'd295/*295:US*/))  xpc10nz <= 9'd296/*296:xpc10nz*/;
                  if ((xpc10nz==9'd296/*296:US*/))  xpc10nz <= 9'd297/*297:xpc10nz*/;
                  if ((xpc10nz==9'd297/*297:US*/))  xpc10nz <= 9'd298/*298:xpc10nz*/;
                  if ((xpc10nz==9'd298/*298:US*/))  xpc10nz <= 9'd299/*299:xpc10nz*/;
                  if ((xpc10nz==9'd299/*299:US*/))  xpc10nz <= 9'd300/*300:xpc10nz*/;
                  if ((xpc10nz==9'd300/*300:US*/))  xpc10nz <= 9'd301/*301:xpc10nz*/;
                  if ((xpc10nz==9'd301/*301:US*/))  xpc10nz <= 9'd302/*302:xpc10nz*/;
                  if ((xpc10nz==9'd302/*302:US*/))  xpc10nz <= 9'd303/*303:xpc10nz*/;
                  if ((xpc10nz==9'd303/*303:US*/))  xpc10nz <= 9'd304/*304:xpc10nz*/;
                  if ((xpc10nz==9'd304/*304:US*/))  xpc10nz <= 9'd305/*305:xpc10nz*/;
                  if ((xpc10nz==9'd305/*305:US*/))  xpc10nz <= 9'd306/*306:xpc10nz*/;
                  if ((xpc10nz==9'd306/*306:US*/))  xpc10nz <= 9'd307/*307:xpc10nz*/;
                  if ((xpc10nz==9'd307/*307:US*/))  xpc10nz <= 9'd308/*308:xpc10nz*/;
                  if ((xpc10nz==9'd308/*308:US*/))  xpc10nz <= 9'd309/*309:xpc10nz*/;
                  if ((xpc10nz==9'd309/*309:US*/))  xpc10nz <= 9'd310/*310:xpc10nz*/;
                  if ((xpc10nz==9'd310/*310:US*/))  xpc10nz <= 9'd311/*311:xpc10nz*/;
                  if ((xpc10nz==9'd311/*311:US*/))  xpc10nz <= 9'd312/*312:xpc10nz*/;
                  if ((xpc10nz==9'd312/*312:US*/))  xpc10nz <= 9'd313/*313:xpc10nz*/;
                  if ((xpc10nz==9'd313/*313:US*/))  xpc10nz <= 9'd314/*314:xpc10nz*/;
                  if ((xpc10nz==9'd314/*314:US*/))  xpc10nz <= 9'd315/*315:xpc10nz*/;
                  if ((xpc10nz==9'd315/*315:US*/))  xpc10nz <= 9'd316/*316:xpc10nz*/;
                  if ((xpc10nz==9'd316/*316:US*/))  xpc10nz <= 9'd317/*317:xpc10nz*/;
                  if ((xpc10nz==9'd317/*317:US*/))  xpc10nz <= 9'd318/*318:xpc10nz*/;
                  if ((xpc10nz==9'd318/*318:US*/))  xpc10nz <= 9'd319/*319:xpc10nz*/;
                  if ((xpc10nz==9'd319/*319:US*/))  xpc10nz <= 9'd320/*320:xpc10nz*/;
                  if ((xpc10nz==9'd320/*320:US*/))  xpc10nz <= 9'd321/*321:xpc10nz*/;
                  if ((xpc10nz==9'd321/*321:US*/))  xpc10nz <= 9'd322/*322:xpc10nz*/;
                  if ((xpc10nz==9'd322/*322:US*/))  xpc10nz <= 9'd323/*323:xpc10nz*/;
                  if ((xpc10nz==9'd323/*323:US*/))  xpc10nz <= 9'd324/*324:xpc10nz*/;
                  if ((xpc10nz==9'd324/*324:US*/))  xpc10nz <= 9'd325/*325:xpc10nz*/;
                  if ((xpc10nz==9'd325/*325:US*/))  xpc10nz <= 9'd326/*326:xpc10nz*/;
                  if ((xpc10nz==9'd326/*326:US*/))  xpc10nz <= 9'd327/*327:xpc10nz*/;
                  if ((xpc10nz==9'd327/*327:US*/))  xpc10nz <= 9'd328/*328:xpc10nz*/;
                  if ((xpc10nz==9'd328/*328:US*/))  xpc10nz <= 9'd329/*329:xpc10nz*/;
                  if ((xpc10nz==9'd329/*329:US*/))  xpc10nz <= 9'd330/*330:xpc10nz*/;
                  if ((xpc10nz==9'd330/*330:US*/))  xpc10nz <= 9'd331/*331:xpc10nz*/;
                  if ((xpc10nz==9'd331/*331:US*/))  xpc10nz <= 9'd332/*332:xpc10nz*/;
                  if ((xpc10nz==9'd332/*332:US*/))  xpc10nz <= 9'd333/*333:xpc10nz*/;
                  if ((xpc10nz==9'd333/*333:US*/))  xpc10nz <= 9'd334/*334:xpc10nz*/;
                  if ((xpc10nz==9'd334/*334:US*/))  xpc10nz <= 9'd335/*335:xpc10nz*/;
                  if ((xpc10nz==9'd335/*335:US*/))  xpc10nz <= 9'd336/*336:xpc10nz*/;
                  if ((xpc10nz==9'd336/*336:US*/))  xpc10nz <= 9'd337/*337:xpc10nz*/;
                  if ((xpc10nz==9'd337/*337:US*/))  xpc10nz <= 9'd338/*338:xpc10nz*/;
                  if ((xpc10nz==9'd338/*338:US*/))  xpc10nz <= 9'd339/*339:xpc10nz*/;
                  if ((xpc10nz==9'd339/*339:US*/))  xpc10nz <= 9'd340/*340:xpc10nz*/;
                  if ((xpc10nz==9'd340/*340:US*/))  xpc10nz <= 9'd341/*341:xpc10nz*/;
                  if ((xpc10nz==9'd341/*341:US*/))  xpc10nz <= 9'd342/*342:xpc10nz*/;
                  if ((xpc10nz==9'd342/*342:US*/))  xpc10nz <= 9'd343/*343:xpc10nz*/;
                  if ((xpc10nz==9'd343/*343:US*/))  xpc10nz <= 9'd344/*344:xpc10nz*/;
                  if ((xpc10nz==9'd344/*344:US*/))  xpc10nz <= 9'd345/*345:xpc10nz*/;
                  if ((xpc10nz==9'd345/*345:US*/))  xpc10nz <= 9'd346/*346:xpc10nz*/;
                  if ((xpc10nz==9'd346/*346:US*/))  xpc10nz <= 9'd347/*347:xpc10nz*/;
                  if ((xpc10nz==9'd347/*347:US*/))  xpc10nz <= 9'd348/*348:xpc10nz*/;
                  if ((xpc10nz==9'd348/*348:US*/))  xpc10nz <= 9'd349/*349:xpc10nz*/;
                  if ((xpc10nz==9'd349/*349:US*/))  xpc10nz <= 9'd350/*350:xpc10nz*/;
                  if ((xpc10nz==9'd350/*350:US*/))  xpc10nz <= 9'd351/*351:xpc10nz*/;
                  if ((xpc10nz==9'd351/*351:US*/))  xpc10nz <= 9'd352/*352:xpc10nz*/;
                  if ((xpc10nz==9'd352/*352:US*/))  xpc10nz <= 9'd353/*353:xpc10nz*/;
                  if ((xpc10nz==9'd353/*353:US*/))  xpc10nz <= 9'd354/*354:xpc10nz*/;
                  if ((xpc10nz==9'd354/*354:US*/))  xpc10nz <= 9'd355/*355:xpc10nz*/;
                  if ((xpc10nz==9'd355/*355:US*/))  xpc10nz <= 9'd356/*356:xpc10nz*/;
                  if ((xpc10nz==9'd356/*356:US*/))  xpc10nz <= 9'd357/*357:xpc10nz*/;
                  if ((xpc10nz==9'd357/*357:US*/))  xpc10nz <= 9'd358/*358:xpc10nz*/;
                  if ((xpc10nz==9'd358/*358:US*/))  xpc10nz <= 9'd359/*359:xpc10nz*/;
                  if ((xpc10nz==9'd359/*359:US*/))  xpc10nz <= 9'd360/*360:xpc10nz*/;
                  if ((xpc10nz==9'd360/*360:US*/))  xpc10nz <= 9'd361/*361:xpc10nz*/;
                  if ((xpc10nz==9'd361/*361:US*/))  xpc10nz <= 9'd362/*362:xpc10nz*/;
                  if ((xpc10nz==9'd362/*362:US*/))  xpc10nz <= 9'd363/*363:xpc10nz*/;
                  if ((xpc10nz==9'd363/*363:US*/))  xpc10nz <= 9'd364/*364:xpc10nz*/;
                  if ((xpc10nz==9'd364/*364:US*/))  xpc10nz <= 9'd365/*365:xpc10nz*/;
                  if ((xpc10nz==9'd365/*365:US*/))  xpc10nz <= 9'd366/*366:xpc10nz*/;
                  if ((xpc10nz==9'd366/*366:US*/))  xpc10nz <= 9'd367/*367:xpc10nz*/;
                  if ((xpc10nz==9'd367/*367:US*/))  xpc10nz <= 9'd368/*368:xpc10nz*/;
                  if ((xpc10nz==9'd368/*368:US*/))  xpc10nz <= 9'd369/*369:xpc10nz*/;
                  if ((xpc10nz==9'd369/*369:US*/))  xpc10nz <= 9'd370/*370:xpc10nz*/;
                  if ((xpc10nz==9'd370/*370:US*/))  xpc10nz <= 9'd371/*371:xpc10nz*/;
                  if ((xpc10nz==9'd371/*371:US*/))  xpc10nz <= 9'd372/*372:xpc10nz*/;
                  if ((xpc10nz==9'd372/*372:US*/))  xpc10nz <= 9'd373/*373:xpc10nz*/;
                  if ((xpc10nz==9'd373/*373:US*/))  xpc10nz <= 9'd374/*374:xpc10nz*/;
                  if ((xpc10nz==9'd374/*374:US*/))  xpc10nz <= 9'd375/*375:xpc10nz*/;
                  if ((xpc10nz==9'd375/*375:US*/))  xpc10nz <= 9'd376/*376:xpc10nz*/;
                  if ((xpc10nz==9'd376/*376:US*/))  xpc10nz <= 9'd377/*377:xpc10nz*/;
                  if ((xpc10nz==9'd377/*377:US*/))  xpc10nz <= 9'd378/*378:xpc10nz*/;
                  if ((xpc10nz==9'd378/*378:US*/))  xpc10nz <= 9'd379/*379:xpc10nz*/;
                  if ((xpc10nz==9'd379/*379:US*/))  xpc10nz <= 9'd380/*380:xpc10nz*/;
                  if ((xpc10nz==9'd380/*380:US*/))  xpc10nz <= 9'd381/*381:xpc10nz*/;
                  if ((xpc10nz==9'd381/*381:US*/))  xpc10nz <= 9'd382/*382:xpc10nz*/;
                  if ((xpc10nz==9'd382/*382:US*/))  xpc10nz <= 9'd383/*383:xpc10nz*/;
                  if ((xpc10nz==9'd383/*383:US*/))  xpc10nz <= 9'd384/*384:xpc10nz*/;
                  if ((xpc10nz==9'd384/*384:US*/))  xpc10nz <= 9'd385/*385:xpc10nz*/;
                  if ((xpc10nz==9'd385/*385:US*/))  xpc10nz <= 9'd386/*386:xpc10nz*/;
                  if ((xpc10nz==9'd386/*386:US*/))  xpc10nz <= 9'd387/*387:xpc10nz*/;
                  if ((xpc10nz==9'd387/*387:US*/))  xpc10nz <= 9'd388/*388:xpc10nz*/;
                  if ((xpc10nz==9'd388/*388:US*/))  xpc10nz <= 9'd389/*389:xpc10nz*/;
                  if ((xpc10nz==9'd389/*389:US*/))  xpc10nz <= 9'd390/*390:xpc10nz*/;
                  if ((xpc10nz==9'd390/*390:US*/))  xpc10nz <= 9'd391/*391:xpc10nz*/;
                  if ((xpc10nz==9'd391/*391:US*/))  xpc10nz <= 9'd392/*392:xpc10nz*/;
                  if ((xpc10nz==9'd392/*392:US*/))  xpc10nz <= 9'd393/*393:xpc10nz*/;
                  if ((xpc10nz==9'd393/*393:US*/))  xpc10nz <= 9'd394/*394:xpc10nz*/;
                  if ((xpc10nz==9'd394/*394:US*/))  xpc10nz <= 9'd395/*395:xpc10nz*/;
                  if ((xpc10nz==9'd395/*395:US*/))  xpc10nz <= 9'd396/*396:xpc10nz*/;
                  if ((xpc10nz==9'd396/*396:US*/))  xpc10nz <= 9'd397/*397:xpc10nz*/;
                  if ((xpc10nz==9'd397/*397:US*/))  xpc10nz <= 9'd398/*398:xpc10nz*/;
                  if ((xpc10nz==9'd398/*398:US*/))  xpc10nz <= 9'd399/*399:xpc10nz*/;
                  if ((xpc10nz==9'd399/*399:US*/))  xpc10nz <= 9'd400/*400:xpc10nz*/;
                  if ((xpc10nz==9'd400/*400:US*/))  xpc10nz <= 9'd497/*497:xpc10nz*/;
                  if ((xpc10nz==9'd402/*402:US*/))  xpc10nz <= 9'd403/*403:xpc10nz*/;
                  if ((xpc10nz==9'd403/*403:US*/))  xpc10nz <= 9'd404/*404:xpc10nz*/;
                  if ((xpc10nz==9'd404/*404:US*/))  xpc10nz <= 9'd405/*405:xpc10nz*/;
                  if ((xpc10nz==9'd406/*406:US*/))  xpc10nz <= 9'd470/*470:xpc10nz*/;
                  if ((xpc10nz==9'd408/*408:US*/))  xpc10nz <= 9'd469/*469:xpc10nz*/;
                  if ((xpc10nz==9'd409/*409:US*/))  xpc10nz <= 9'd410/*410:xpc10nz*/;
                  if ((xpc10nz==9'd411/*411:US*/))  xpc10nz <= 9'd412/*412:xpc10nz*/;
                  if ((xpc10nz==9'd412/*412:US*/))  xpc10nz <= 9'd413/*413:xpc10nz*/;
                  if ((xpc10nz==9'd413/*413:US*/))  xpc10nz <= 9'd414/*414:xpc10nz*/;
                  if ((xpc10nz==9'd415/*415:US*/))  xpc10nz <= 9'd465/*465:xpc10nz*/;
                  if ((xpc10nz==9'd416/*416:US*/))  xpc10nz <= 9'd417/*417:xpc10nz*/;
                  if ((xpc10nz==9'd417/*417:US*/))  xpc10nz <= 9'd418/*418:xpc10nz*/;
                  if ((xpc10nz==9'd418/*418:US*/))  xpc10nz <= 9'd419/*419:xpc10nz*/;
                  if ((xpc10nz==9'd420/*420:US*/))  xpc10nz <= 9'd411/*411:xpc10nz*/;
                  if ((xpc10nz==9'd421/*421:US*/))  xpc10nz <= 9'd411/*411:xpc10nz*/;
                  if ((xpc10nz==9'd422/*422:US*/))  xpc10nz <= 9'd423/*423:xpc10nz*/;
                  if ((xpc10nz==9'd423/*423:US*/))  xpc10nz <= 9'd424/*424:xpc10nz*/;
                  if ((xpc10nz==9'd424/*424:US*/))  xpc10nz <= 9'd425/*425:xpc10nz*/;
                  if ((xpc10nz==9'd426/*426:US*/))  xpc10nz <= 9'd427/*427:xpc10nz*/;
                  if ((xpc10nz==9'd427/*427:US*/))  xpc10nz <= 9'd428/*428:xpc10nz*/;
                  if ((xpc10nz==9'd428/*428:US*/))  xpc10nz <= 9'd429/*429:xpc10nz*/;
                  if ((xpc10nz==9'd430/*430:US*/))  xpc10nz <= 9'd431/*431:xpc10nz*/;
                  if ((xpc10nz==9'd431/*431:US*/))  xpc10nz <= 9'd432/*432:xpc10nz*/;
                  if ((xpc10nz==9'd432/*432:US*/))  xpc10nz <= 9'd433/*433:xpc10nz*/;
                  if ((xpc10nz==9'd434/*434:US*/))  xpc10nz <= 9'd426/*426:xpc10nz*/;
                  if ((xpc10nz==9'd435/*435:US*/))  xpc10nz <= 9'd426/*426:xpc10nz*/;
                  if ((xpc10nz==9'd436/*436:US*/))  xpc10nz <= 9'd437/*437:xpc10nz*/;
                  if ((xpc10nz==9'd437/*437:US*/))  xpc10nz <= 9'd438/*438:xpc10nz*/;
                  if ((xpc10nz==9'd438/*438:US*/))  xpc10nz <= 9'd439/*439:xpc10nz*/;
                  if ((xpc10nz==9'd440/*440:US*/))  xpc10nz <= 9'd430/*430:xpc10nz*/;
                  if ((xpc10nz==9'd441/*441:US*/))  xpc10nz <= 9'd430/*430:xpc10nz*/;
                  if ((xpc10nz==9'd442/*442:US*/))  xpc10nz <= 9'd443/*443:xpc10nz*/;
                  if ((xpc10nz==9'd443/*443:US*/))  xpc10nz <= 9'd444/*444:xpc10nz*/;
                  if ((xpc10nz==9'd444/*444:US*/))  xpc10nz <= 9'd445/*445:xpc10nz*/;
                  if ((xpc10nz==9'd447/*447:US*/))  xpc10nz <= 9'd448/*448:xpc10nz*/;
                  if ((xpc10nz==9'd450/*450:US*/))  xpc10nz <= 9'd451/*451:xpc10nz*/;
                  if ((xpc10nz==9'd453/*453:US*/))  xpc10nz <= 9'd454/*454:xpc10nz*/;
                  if ((xpc10nz==9'd456/*456:US*/))  xpc10nz <= 9'd457/*457:xpc10nz*/;
                  if ((xpc10nz==9'd460/*460:US*/))  xpc10nz <= 9'd461/*461:xpc10nz*/;
                  if ((xpc10nz==9'd461/*461:US*/))  xpc10nz <= 9'd462/*462:xpc10nz*/;
                  if ((xpc10nz==9'd473/*473:US*/))  xpc10nz <= 9'd474/*474:xpc10nz*/;
                  if ((xpc10nz==9'd477/*477:US*/))  xpc10nz <= 9'd478/*478:xpc10nz*/;
                  if ((xpc10nz==9'd481/*481:US*/))  xpc10nz <= 9'd482/*482:xpc10nz*/;
                  if ((xpc10nz==9'd484/*484:US*/))  xpc10nz <= 9'd485/*485:xpc10nz*/;
                  if ((xpc10nz==9'd487/*487:US*/))  xpc10nz <= 9'd488/*488:xpc10nz*/;
                  if ((xpc10nz==9'd490/*490:US*/))  xpc10nz <= 9'd489/*489:xpc10nz*/;
                  if ((xpc10nz==9'd493/*493:US*/))  xpc10nz <= 9'd491/*491:xpc10nz*/;
                  if ((xpc10nz==9'd494/*494:US*/))  xpc10nz <= 9'd401/*401:xpc10nz*/;
                  if ((xpc10nz==9'd495/*495:US*/))  xpc10nz <= 9'd496/*496:xpc10nz*/;
                  if ((xpc10nz==9'd497/*497:US*/))  xpc10nz <= 9'd495/*495:xpc10nz*/;
                   end 
              //End structure HPR sw_test.exe


       end 
      

  CV_SP_SSRAM_FL1 #(6'd32, 4'd9, 9'd510, 6'd32) A_UINT_CC_SCALbx34_ARA0(clk, reset, A_UINT_CC_SCALbx34_ARA0_RDD0, A_UINT_CC_SCALbx34_ARA0_AD0
, A_UINT_CC_SCALbx34_ARA0_WEN0, A_UINT_CC_SCALbx34_ARA0_REN0, A_UINT_CC_SCALbx34_ARA0_WRD0);

  CV_SP_SSRAM_FL1 #(6'd32, 4'd10, 10'd798, 6'd32) A_SINT_CC_SCALbx16_ARA0(clk, reset, A_SINT_CC_SCALbx16_ARA0_RDD0, A_SINT_CC_SCALbx16_ARA0_AD0
, A_SINT_CC_SCALbx16_ARA0_WEN0, A_SINT_CC_SCALbx16_ARA0_REN0, A_SINT_CC_SCALbx16_ARA0_WRD0);

  CV_SP_SSRAM_FL1 #(5'd16, 4'd8, 8'd148, 5'd16) A_16_SS_CC_SCALbx10_ARA0(clk, reset, A_16_SS_CC_SCALbx10_ARA0_RDD0, A_16_SS_CC_SCALbx10_ARA0_AD0
, A_16_SS_CC_SCALbx10_ARA0_WEN0, A_16_SS_CC_SCALbx10_ARA0_REN0, A_16_SS_CC_SCALbx10_ARA0_WRD0);

  CV_SP_SSRAM_FL1 #(5'd16, 4'd8, 8'd152, 5'd16) A_16_SS_CC_SCALbx14_ARC0(clk, reset, A_16_SS_CC_SCALbx14_ARC0_RDD0, A_16_SS_CC_SCALbx14_ARC0_AD0
, A_16_SS_CC_SCALbx14_ARC0_WEN0, A_16_SS_CC_SCALbx14_ARC0_REN0, A_16_SS_CC_SCALbx14_ARC0_WRD0);

  CV_SP_SSRAM_FL1 #(5'd16, 3'd6, 6'd38, 5'd16) A_16_SS_CC_SCALbx12_ARB0(clk, reset, A_16_SS_CC_SCALbx12_ARB0_RDD0, A_16_SS_CC_SCALbx12_ARB0_AD0
, A_16_SS_CC_SCALbx12_ARB0_WEN0, A_16_SS_CC_SCALbx12_ARB0_REN0, A_16_SS_CC_SCALbx12_ARB0_WRD0);

  CV_INT_FL2_MULTIPLIER_US i302CV_INT_FL2_MULTIPLIER_US(clk, reset, iuMULTIPLIER10_RR, iuMULTIPLIER10_NN, iuMULTIPLIER10_DD, iuMULTIPLIER10_err
);
  CV_SP_SSRAM_FL1 #(7'd64, 4'd8, 8'd156, 7'd64) A_64_SS_CC_SCALbx52_ARA0(clk, reset, A_64_SS_CC_SCALbx52_ARA0_RDD0, A_64_SS_CC_SCALbx52_ARA0_AD0
, A_64_SS_CC_SCALbx52_ARA0_WEN0, A_64_SS_CC_SCALbx52_ARA0_REN0, A_64_SS_CC_SCALbx52_ARA0_WRD0);

  CV_INT_FL2_MULTIPLIER_US i300CV_INT_FL2_MULTIPLIER_US(clk, reset, iuMULTIPLIER12_RR, iuMULTIPLIER12_NN, iuMULTIPLIER12_DD, iuMULTIPLIER12_err
);
  CV_SP_SSRAM_FL1 #(7'd64, 4'd8, 8'd156, 7'd64) A_64_SS_CC_SCALbx54_ARB0(clk, reset, A_64_SS_CC_SCALbx54_ARB0_RDD0, A_64_SS_CC_SCALbx54_ARB0_AD0
, A_64_SS_CC_SCALbx54_ARB0_WEN0, A_64_SS_CC_SCALbx54_ARB0_REN0, A_64_SS_CC_SCALbx54_ARB0_WRD0);

  CV_INT_FL2_MULTIPLIER_US i298CV_INT_FL2_MULTIPLIER_US(clk, reset, iuMULTIPLIER14_RR, iuMULTIPLIER14_NN, iuMULTIPLIER14_DD, iuMULTIPLIER14_err
);
  CV_SP_SSRAM_FL1 #(7'd64, 4'd8, 8'd156, 7'd64) A_64_SS_CC_SCALbx56_ARC0(clk, reset, A_64_SS_CC_SCALbx56_ARC0_RDD0, A_64_SS_CC_SCALbx56_ARC0_AD0
, A_64_SS_CC_SCALbx56_ARC0_WEN0, A_64_SS_CC_SCALbx56_ARC0_REN0, A_64_SS_CC_SCALbx56_ARC0_WRD0);

  CV_SP_SSRAM_FL1 #(7'd64, 4'd8, 8'd156, 7'd64) A_64_SS_CC_SCALbx58_ARD0(clk, reset, A_64_SS_CC_SCALbx58_ARD0_RDD0, A_64_SS_CC_SCALbx58_ARD0_AD0
, A_64_SS_CC_SCALbx58_ARD0_WEN0, A_64_SS_CC_SCALbx58_ARD0_REN0, A_64_SS_CC_SCALbx58_ARD0_WRD0);

  CV_SP_SSRAM_FL1 #(6'd32, 3'd7, 7'd77, 6'd32) A_SINT_CC_SCALbx26_ARJ0(clk, reset, A_SINT_CC_SCALbx26_ARJ0_RDD0, A_SINT_CC_SCALbx26_ARJ0_AD0
, A_SINT_CC_SCALbx26_ARJ0_WEN0, A_SINT_CC_SCALbx26_ARJ0_REN0, A_SINT_CC_SCALbx26_ARJ0_WRD0);

always @(*) xpc10_stall = ((xpc10nz==9'd449/*449:US*/) || (xpc10nz==9'd451/*451:US*/) || (xpc10nz==9'd454/*454:US*/) || (xpc10nz==9'd457/*457:US*/) || (xpc10nz
==9'd474/*474:US*/) || (xpc10nz==9'd478/*478:US*/) || (xpc10nz==9'd482/*482:US*/) || (xpc10nz==9'd485/*485:US*/) || (xpc10nz==9'd488/*488:US*/)) && 
!UINTCCSCALbx34ARA0RRh12shot0 || ((xpc10nz==9'd448/*448:US*/) || (xpc10nz==9'd452/*452:US*/) || (xpc10nz==9'd455/*455:US*/) || (xpc10nz
==9'd458/*458:US*/) || (xpc10nz==9'd475/*475:US*/) || (xpc10nz==9'd479/*479:US*/) || (xpc10nz==9'd483/*483:US*/)) && !UINTCCSCALbx34ARA0RRh10shot0
 || ((xpc10nz==9'd414/*414:US*/) || (xpc10nz==9'd425/*425:US*/) || (xpc10nz==9'd445/*445:US*/) || (xpc10nz==9'd462/*462:US*/)) && !Z64SSCCSCALbx54ARB0RRh10shot0
 || ((xpc10nz==9'd496/*496:US*/) || (xpc10nz==9'd410/*410:US*/)) && !Z16SSCCSCALbx12ARB0RRh10shot0 || ((xpc10nz==9'd433/*433:US*/) || 
(xpc10nz==9'd429/*429:US*/)) && !Z64SSCCSCALbx56ARC0RRh10shot0 || ((xpc10nz==9'd439/*439:US*/) || (xpc10nz==9'd429/*429:US*/)) && !Z64SSCCSCALbx58ARD0RRh10shot0
 || ((xpc10nz==9'd439/*439:US*/) || (xpc10nz==9'd433/*433:US*/)) && !Z64SSCCSCALbx52ARA0RRh10shot0 || !SINTCCSCALbx16ARA0RRh10shot0 && 
(xpc10nz==9'd419/*419:US*/) || !Z16SSCCSCALbx14ARC0RRh10shot0 && (xpc10nz==9'd496/*496:US*/) || !Z16SSCCSCALbx10ARA0RRh10shot0 && (xpc10nz
==9'd410/*410:US*/);

// 2 vectors of width 9
// 38 vectors of width 1
// 25 vectors of width 32
// 6 vectors of width 16
// 10 vectors of width 64
// 1 vectors of width 7
// 12 vectors of width 8
// 1 vectors of width 6
// 1 vectors of width 10
// 608 bits in scalar variables
// Total state bits in module = 2319 bits.
// 501 continuously assigned (wire/non-state) bits 
//   cell CV_SP_SSRAM_FL1 count=10
//   cell CV_INT_FL2_MULTIPLIER_US count=3
// Total number of leaf cells = 2
endmodule

// 
/*

// Highest off-chip SRAM/DRAM location in use on port dram0bank is <null> (--not-used--) bytes=1048576
// res3: Thread=xpc10 state=X1:"1:xpc10:1"
*-----+-----+---------+-------*
| npc | eno | Phaser  | Work  |
*-----+-----+---------+-------*
| 497 | -   | R0 CTRL |       |
| 497 | 959 | R0 DATA |       |
| 497 | 959 | W0 DATA | EXEC  |
*-----+-----+---------+-------*

// res3: Thread=xpc10 state=X2:"2:xpc10:2"
*-----+-----+---------+---------------------------------------------------------------------------------------------------------------------------------*
| npc | eno | Phaser  | Work                                                                                                                            |
*-----+-----+---------+---------------------------------------------------------------------------------------------------------------------------------*
| 495 | -   | R0 CTRL | @16_SS/CC/SCALbx14_ARC0 te=495-te-495 read args=0, TSPin0.6_V_0;@16_SS/CC/SCALbx12_ARB0 te=495-te-495 read args=0, TSPen1.8_V_0 |
| 496 | -   | R1 CTRL |                                                                                                                                 |
| 496 | 957 | R1 DATA |                                                                                                                                 |
| 496 | 957 | W0 DATA | EXEC ;TSPe1._SPILL_256 te=496-te-496 scalarw args=C(TSPen1.8_V_0)                                                               |
| 496 | 958 | R1 DATA |                                                                                                                                 |
| 496 | 958 | W0 DATA | EXEC ;TSPen1.8_V_0 te=496-te-496 scalarw args=C(1+TSPen1.8_V_0)                                                                 |
*-----+-----+---------+---------------------------------------------------------------------------------------------------------------------------------*

// res3: Thread=xpc10 state=X3:"3:xpc10:3"
*-----+-----+---------+--------------------------------------------------------------------------------------------------------------------------------------------------------------------------*
| npc | eno | Phaser  | Work                                                                                                                                                                     |
*-----+-----+---------+--------------------------------------------------------------------------------------------------------------------------------------------------------------------------*
| 492 | -   | R0 CTRL |                                                                                                                                                                          |
| 492 | 955 | R0 DATA |                                                                                                                                                                          |
| 492 | 955 | W0 DATA | EXEC ;TSPin0.6_V_0 te=492-te-492 scalarw args=C(1+TSPin0.6_V_0);phase te=492-te-492 scalarw args=Cu(3);@_SINT/CC/SCALbx26_ARJ0 te=492-te-492 write args=0, TSPin0.6_V_0\ |
|     |     |         | , C(TSPe1._SPILL_256);TSPru0.12_V_0 te=492-te-492 scalarw args=C(0) W/P:waypoint %u %u                                                                                   |
| 493 | 955 | W1 DATA |                                                                                                                                                                          |
| 492 | 956 | R0 DATA |                                                                                                                                                                          |
| 492 | 956 | W0 DATA | EXEC ;TSPen1.8_V_0 te=492-te-492 scalarw args=C(0);TSPin0.6_V_0 te=492-te-492 scalarw args=C(1+TSPin0.6_V_0);@_SINT/CC/SCALbx26_ARJ0 te=492-te-492 write args=0, TSPin0\ |
|     |     |         | .6_V_0, C(TSPe1._SPILL_256)                                                                                                                                              |
| 494 | 956 | W1 DATA |                                                                                                                                                                          |
*-----+-----+---------+--------------------------------------------------------------------------------------------------------------------------------------------------------------------------*

// res3: Thread=xpc10 state=X4:"4:xpc10:4"
*-----+-----+---------+-------------------------------------------------------------------------------------------------------------------------------------*
| npc | eno | Phaser  | Work                                                                                                                                |
*-----+-----+---------+-------------------------------------------------------------------------------------------------------------------------------------*
| 491 | -   | R0 CTRL |                                                                                                                                     |
| 491 | 953 | R0 DATA |                                                                                                                                     |
| 491 | 953 | W0 DATA | EXEC ;phase te=491-te-491 scalarw args=Cu(12);@_UINT/CC/SCALbx38_crc_reg te=491-te-491 scalarw args=Cu(-1) W/P:crc reg now:  reg=%H |
| 491 | 954 | R0 DATA |                                                                                                                                     |
| 491 | 954 | W0 DATA | EXEC                                                                                                                                |
*-----+-----+---------+-------------------------------------------------------------------------------------------------------------------------------------*

// res3: Thread=xpc10 state=X5:"5:xpc10:5"
*-----+-----+---------+-------*
| npc | eno | Phaser  | Work  |
*-----+-----+---------+-------*
| 490 | -   | R0 CTRL |       |
| 490 | 952 | R0 DATA |       |
| 490 | 952 | W0 DATA | EXEC  |
*-----+-----+---------+-------*

// res3: Thread=xpc10 state=X6:"6:xpc10:6"
*-----+-----+---------+--------------------------------------------------------------------*
| npc | eno | Phaser  | Work                                                               |
*-----+-----+---------+--------------------------------------------------------------------*
| 489 | -   | R0 CTRL |                                                                    |
| 489 | 951 | R0 DATA |                                                                    |
| 489 | 951 | W0 DATA | EXEC ;@_UINT/CC/SCALbx38_crc_reg te=489-te-489 scalarw args=Cu(-1) |
*-----+-----+---------+--------------------------------------------------------------------*

// res3: Thread=xpc10 state=X7:"7:xpc10:7"
*-----+-----+---------+--------------------------------------------------------*
| npc | eno | Phaser  | Work                                                   |
*-----+-----+---------+--------------------------------------------------------*
| 487 | -   | R0 CTRL |                                                        |
| 487 | 950 | R0 DATA | @_UINT/CC/SCALbx34_ARA0 te=487-te-487 read args=0, 255 |
| 488 | 950 | R1 DATA |                                                        |
| 488 | 950 | W0 DATA | EXEC  W/P:self test startup %d...                      |
*-----+-----+---------+--------------------------------------------------------*

// res3: Thread=xpc10 state=X8:"8:xpc10:8"
*-----+-----+---------+-----------------------------------*
| npc | eno | Phaser  | Work                              |
*-----+-----+---------+-----------------------------------*
| 486 | -   | R0 CTRL |                                   |
| 486 | 949 | R0 DATA |                                   |
| 486 | 949 | W0 DATA | EXEC  W/P:self test startup %d... |
*-----+-----+---------+-----------------------------------*

// res3: Thread=xpc10 state=X9:"9:xpc10:9"
*-----+-----+---------+--------------------------------------------------------------------------------------------*
| npc | eno | Phaser  | Work                                                                                       |
*-----+-----+---------+--------------------------------------------------------------------------------------------*
| 484 | -   | R0 CTRL |                                                                                            |
| 484 | 948 | R0 DATA | @_UINT/CC/SCALbx34_ARA0 te=484-te-484 read args=0, 255                                     |
| 485 | 948 | R1 DATA |                                                                                            |
| 485 | 948 | W0 DATA | EXEC ;@_UINT/CC/SCALbx38_byteno te=485-te-485 scalarw args=E54 W/P:self test startup %d... |
*-----+-----+---------+--------------------------------------------------------------------------------------------*

// res3: Thread=xpc10 state=X10:"10:xpc10:10"
*-----+-----+---------+---------------------------------------------------------------------------------------------*
| npc | eno | Phaser  | Work                                                                                        |
*-----+-----+---------+---------------------------------------------------------------------------------------------*
| 481 | -   | R0 CTRL |                                                                                             |
| 481 | 947 | R0 DATA | @_UINT/CC/SCALbx34_ARA0 te=481-te-481 read args=0, 1                                        |
| 482 | 947 | R1 DATA | @_UINT/CC/SCALbx34_ARA0 te=482-te-482 read args=0, 255                                      |
| 483 | 947 | R2 DATA |                                                                                             |
| 483 | 947 | W0 DATA | EXEC ;@_UINT/CC/SCALbx38_crc_reg te=483-te-483 scalarw args=E57 W/P:crc update hex:  reg... |
*-----+-----+---------+---------------------------------------------------------------------------------------------*

// res3: Thread=xpc10 state=X11:"11:xpc10:11"
*-----+-----+---------+------------------------------------------------------------------------------------------------------------*
| npc | eno | Phaser  | Work                                                                                                       |
*-----+-----+---------+------------------------------------------------------------------------------------------------------------*
| 480 | -   | R0 CTRL |                                                                                                            |
| 480 | 946 | R0 DATA |                                                                                                            |
| 480 | 946 | W0 DATA | EXEC ;@_UINT/CC/SCALbx38_byteno te=480-te-480 scalarw args=E54;TCpr0.40_V_0 te=480-te-480 scalarw args=E55 |
*-----+-----+---------+------------------------------------------------------------------------------------------------------------*

// res3: Thread=xpc10 state=X12:"12:xpc10:12"
*-----+-----+---------+---------------------------------------------------------------------------------------------*
| npc | eno | Phaser  | Work                                                                                        |
*-----+-----+---------+---------------------------------------------------------------------------------------------*
| 477 | -   | R0 CTRL |                                                                                             |
| 477 | 945 | R0 DATA | @_UINT/CC/SCALbx34_ARA0 te=477-te-477 read args=0, 128                                      |
| 478 | 945 | R1 DATA | @_UINT/CC/SCALbx34_ARA0 te=478-te-478 read args=0, TCpr0.40_V_0                             |
| 479 | 945 | R2 DATA |                                                                                             |
| 479 | 945 | W0 DATA | EXEC ;@_UINT/CC/SCALbx38_crc_reg te=479-te-479 scalarw args=E56 W/P:crc update hex:  reg... |
*-----+-----+---------+---------------------------------------------------------------------------------------------*

// res3: Thread=xpc10 state=X13:"13:xpc10:13"
*-----+-----+---------+------------------------------------------------------------------------------------------------------------*
| npc | eno | Phaser  | Work                                                                                                       |
*-----+-----+---------+------------------------------------------------------------------------------------------------------------*
| 476 | -   | R0 CTRL |                                                                                                            |
| 476 | 944 | R0 DATA |                                                                                                            |
| 476 | 944 | W0 DATA | EXEC ;@_UINT/CC/SCALbx38_byteno te=476-te-476 scalarw args=E54;TCpr0.44_V_0 te=476-te-476 scalarw args=E55 |
*-----+-----+---------+------------------------------------------------------------------------------------------------------------*

// res3: Thread=xpc10 state=X14:"14:xpc10:14"
*-----+-----+---------+---------------------------------------------------------------------------------------------*
| npc | eno | Phaser  | Work                                                                                        |
*-----+-----+---------+---------------------------------------------------------------------------------------------*
| 473 | -   | R0 CTRL |                                                                                             |
| 473 | 943 | R0 DATA | @_UINT/CC/SCALbx34_ARA0 te=473-te-473 read args=0, 1                                        |
| 474 | 943 | R1 DATA | @_UINT/CC/SCALbx34_ARA0 te=474-te-474 read args=0, TCpr0.44_V_0                             |
| 475 | 943 | R2 DATA |                                                                                             |
| 475 | 943 | W0 DATA | EXEC ;@_UINT/CC/SCALbx38_crc_reg te=475-te-475 scalarw args=E53 W/P:crc update hex:  reg... |
*-----+-----+---------+---------------------------------------------------------------------------------------------*

// res3: Thread=xpc10 state=X15:"15:xpc10:15"
*-----+-----+---------+------------------------------*
| npc | eno | Phaser  | Work                         |
*-----+-----+---------+------------------------------*
| 472 | -   | R0 CTRL |                              |
| 472 | 942 | R0 DATA |                              |
| 472 | 942 | W0 DATA | EXEC  W/P:GSAI:hpr_sysexit:0 |
*-----+-----+---------+------------------------------*

// res3: Thread=xpc10 state=X16:"16:xpc10:16"
*-----+-----+---------+----------------------------------------------------*
| npc | eno | Phaser  | Work                                               |
*-----+-----+---------+----------------------------------------------------*
| 471 | -   | R0 CTRL |                                                    |
| 471 | 941 | R0 DATA |                                                    |
| 471 | 941 | W0 DATA | EXEC ;TSPsw1.2_V_0 te=471-te-471 scalarw args=C(0) |
*-----+-----+---------+----------------------------------------------------*

// res3: Thread=xpc10 state=X17:"17:xpc10:17"
*-----+-----+---------+----------------------------------------------------*
| npc | eno | Phaser  | Work                                               |
*-----+-----+---------+----------------------------------------------------*
| 470 | -   | R0 CTRL |                                                    |
| 470 | 939 | R0 DATA |                                                    |
| 470 | 939 | W0 DATA | EXEC ;TSPsw1.2_V_1 te=470-te-470 scalarw args=C(1) |
| 470 | 940 | R0 DATA |                                                    |
| 470 | 940 | W0 DATA | EXEC                                               |
*-----+-----+---------+----------------------------------------------------*

// res3: Thread=xpc10 state=X18:"18:xpc10:18"
*-----+-----+---------+-----------------------------------------------------*
| npc | eno | Phaser  | Work                                                |
*-----+-----+---------+-----------------------------------------------------*
| 469 | -   | R0 CTRL |                                                     |
| 469 | 937 | R0 DATA |                                                     |
| 469 | 937 | W0 DATA | EXEC ;TSPru0.12_V_1 te=469-te-469 scalarw args=C(0) |
| 469 | 938 | R0 DATA |                                                     |
| 469 | 938 | W0 DATA | EXEC                                                |
*-----+-----+---------+-----------------------------------------------------*

// res3: Thread=xpc10 state=X19:"19:xpc10:19"
*-----+-----+---------+-------------------------------------------------------------------------------------------------------------------------------------------------------------*
| npc | eno | Phaser  | Work                                                                                                                                                        |
*-----+-----+---------+-------------------------------------------------------------------------------------------------------------------------------------------------------------*
| 468 | -   | R0 CTRL |                                                                                                                                                             |
| 468 | 935 | R0 DATA |                                                                                                                                                             |
| 468 | 935 | W0 DATA | EXEC ;TSPru0.12_V_0 te=468-te-468 scalarw args=C(1+TSPru0.12_V_0)                                                                                           |
| 468 | 936 | R0 DATA |                                                                                                                                                             |
| 468 | 936 | W0 DATA | EXEC ;phase te=468-te-468 scalarw args=Cu(4);TSPen0.17_V_0 te=468-te-468 scalarw args=C(0);TSPne2.10_V_1 te=468-te-468 scalarw args=C((1+TSPru0.12_V_1)%2)\ |
|     |     |         | ;TSPne2.10_V_0 te=468-te-468 scalarw args=C(TSPru0.12_V_1%2) W/P:waypoint %u %u                                                                             |
*-----+-----+---------+-------------------------------------------------------------------------------------------------------------------------------------------------------------*

// res3: Thread=xpc10 state=X20:"20:xpc10:20"
*-----+-----+---------+--------------------------------------------------------*
| npc | eno | Phaser  | Work                                                   |
*-----+-----+---------+--------------------------------------------------------*
| 467 | -   | R0 CTRL |                                                        |
| 467 | 933 | R0 DATA |                                                        |
| 467 | 933 | W0 DATA | EXEC ;TSPe0._SPILL_256 te=467-te-467 scalarw args=C(0) |
| 467 | 934 | R0 DATA |                                                        |
| 467 | 934 | W0 DATA | EXEC                                                   |
*-----+-----+---------+--------------------------------------------------------*

// res3: Thread=xpc10 state=X21:"21:xpc10:21"
*-----+-----+---------+------------------------------------------------------------------------------------------------------------------*
| npc | eno | Phaser  | Work                                                                                                             |
*-----+-----+---------+------------------------------------------------------------------------------------------------------------------*
| 466 | -   | R0 CTRL |                                                                                                                  |
| 466 | 932 | R0 DATA |                                                                                                                  |
| 466 | 932 | W0 DATA | EXEC ;TSPne2.10_V_3 te=466-te-466 scalarw args=C(0);TSPne2.10_V_2 te=466-te-466 scalarw args=C(TSPe0._SPILL_256) |
*-----+-----+---------+------------------------------------------------------------------------------------------------------------------*

// res3: Thread=xpc10 state=X22:"22:xpc10:22"
*-----+-----+---------+-------------------------------------------------------------------------------------------------------------------------------------*
| npc | eno | Phaser  | Work                                                                                                                                |
*-----+-----+---------+-------------------------------------------------------------------------------------------------------------------------------------*
| 465 | -   | R0 CTRL |                                                                                                                                     |
| 465 | 930 | R0 DATA |                                                                                                                                     |
| 465 | 930 | W0 DATA | EXEC ;phase te=465-te-465 scalarw args=Cu(8+256*TSPru0.12_V_1);TSPte2.13_V_0 te=465-te-465 scalarw args=C(0) W/P:Scored h matrix %u |
| 465 | 931 | R0 DATA |                                                                                                                                     |
| 465 | 931 | W0 DATA | EXEC                                                                                                                                |
*-----+-----+---------+-------------------------------------------------------------------------------------------------------------------------------------*

// res3: Thread=xpc10 state=X23:"23:xpc10:23"
*-----+-----+---------+-------------------------------------------------------------------------------------------------------------------------------------------------------*
| npc | eno | Phaser  | Work                                                                                                                                                  |
*-----+-----+---------+-------------------------------------------------------------------------------------------------------------------------------------------------------*
| 464 | -   | R0 CTRL |                                                                                                                                                       |
| 464 | 928 | R0 DATA |                                                                                                                                                       |
| 464 | 928 | W0 DATA | EXEC ;phase te=464-te-464 scalarw args=Cu(10+256*TSPru0.12_V_1);@_UINT/CC/SCALbx36_crc_reg te=464-te-464 scalarw args=Cu(-1) W/P:crc reg now:  reg=%H |
| 464 | 929 | R0 DATA |                                                                                                                                                       |
| 464 | 929 | W0 DATA | EXEC ;TSPte2.13_V_2 te=464-te-464 scalarw args=C(0);TSPte2.13_V_1 te=464-te-464 scalarw args=E52                                                      |
*-----+-----+---------+-------------------------------------------------------------------------------------------------------------------------------------------------------*

// res3: Thread=xpc10 state=X24:"24:xpc10:24"
*-----+-----+---------+---------------------------------------------------------------------------------------------------------------------*
| npc | eno | Phaser  | Work                                                                                                                |
*-----+-----+---------+---------------------------------------------------------------------------------------------------------------------*
| 463 | -   | R0 CTRL |                                                                                                                     |
| 463 | 927 | R0 DATA |                                                                                                                     |
| 463 | 927 | W0 DATA | EXEC ;TSPcr2.16_V_1 te=463-te-463 scalarw args=C(0);TSPcr2.16_V_0 te=463-te-463 scalarw args=C((1+TSPru0.12_V_1)%2) |
*-----+-----+---------+---------------------------------------------------------------------------------------------------------------------*

// res3: Thread=xpc10 state=X25:"25:xpc10:25"
*-----+-----+---------+-------------------------------------------------------------------------------------------------------------------------*
| npc | eno | Phaser  | Work                                                                                                                    |
*-----+-----+---------+-------------------------------------------------------------------------------------------------------------------------*
| 459 | -   | R0 CTRL |                                                                                                                         |
| 459 | 925 | R0 DATA |                                                                                                                         |
| 459 | 925 | W0 DATA | EXEC ;d_monitor te=459-te-459 scalarw args=E48;TSPru0.12_V_1 te=459-te-459 scalarw args=C(1+TSPru0.12_V_1) W/P:step %u\ |
|     |     |         |  crc is %d   ...                                                                                                        |
| 459 | 926 | R0 DATA | iuMULTIPLIER14 te=459-te-459 *fixed-function-structural-alu* args=C64u(TSPcr2.16_V_0), E2                               |
| 460 | 926 | R1 DATA |                                                                                                                         |
| 461 | 926 | R2 DATA | @64_SS/CC/SCALbx54_ARB0 te=461-te-461 read args=0, E49                                                                  |
| 462 | 926 | R3 DATA |                                                                                                                         |
| 462 | 926 | W0 DATA | EXEC ;@_UINT/CC/SCALbx36_byteno te=462-te-462 scalarw args=E41;TCpr0.13_V_0 te=462-te-462 scalarw args=E50;TSPcr2.16_V\ |
|     |     |         | _2 te=462-te-462 scalarw args=E51 W/P:process unit word %d...                                                           |
*-----+-----+---------+-------------------------------------------------------------------------------------------------------------------------*

// res3: Thread=xpc10 state=X26:"26:xpc10:26"
*-----+-----+---------+----------------------------------------------------------------------------------------------------------------------------------*
| npc | eno | Phaser  | Work                                                                                                                             |
*-----+-----+---------+----------------------------------------------------------------------------------------------------------------------------------*
| 456 | -   | R0 CTRL |                                                                                                                                  |
| 456 | 924 | R0 DATA | @_UINT/CC/SCALbx34_ARA0 te=456-te-456 read args=0, E37                                                                           |
| 457 | 924 | R1 DATA | @_UINT/CC/SCALbx34_ARA0 te=457-te-457 read args=0, TCpr0.13_V_0                                                                  |
| 458 | 924 | R2 DATA |                                                                                                                                  |
| 458 | 924 | W0 DATA | EXEC ;@_UINT/CC/SCALbx36_crc_reg te=458-te-458 scalarw args=E46;@_UINT/CC/SCALbx36_byteno te=458-te-458 scalarw args=E41;TCpr0.\ |
|     |     |         | 21_V_0 te=458-te-458 scalarw args=E47 W/P:crc update hex:  reg...                                                                |
*-----+-----+---------+----------------------------------------------------------------------------------------------------------------------------------*

// res3: Thread=xpc10 state=X27:"27:xpc10:27"
*-----+-----+---------+----------------------------------------------------------------------------------------------------------------------------------*
| npc | eno | Phaser  | Work                                                                                                                             |
*-----+-----+---------+----------------------------------------------------------------------------------------------------------------------------------*
| 453 | -   | R0 CTRL |                                                                                                                                  |
| 453 | 923 | R0 DATA | @_UINT/CC/SCALbx34_ARA0 te=453-te-453 read args=0, E43                                                                           |
| 454 | 923 | R1 DATA | @_UINT/CC/SCALbx34_ARA0 te=454-te-454 read args=0, TCpr0.21_V_0                                                                  |
| 455 | 923 | R2 DATA |                                                                                                                                  |
| 455 | 923 | W0 DATA | EXEC ;@_UINT/CC/SCALbx36_crc_reg te=455-te-455 scalarw args=E44;@_UINT/CC/SCALbx36_byteno te=455-te-455 scalarw args=E41;TCpr0.\ |
|     |     |         | 29_V_0 te=455-te-455 scalarw args=E45 W/P:crc update hex:  reg...                                                                |
*-----+-----+---------+----------------------------------------------------------------------------------------------------------------------------------*

// res3: Thread=xpc10 state=X28:"28:xpc10:28"
*-----+-----+---------+----------------------------------------------------------------------------------------------------------------------------------*
| npc | eno | Phaser  | Work                                                                                                                             |
*-----+-----+---------+----------------------------------------------------------------------------------------------------------------------------------*
| 450 | -   | R0 CTRL |                                                                                                                                  |
| 450 | 922 | R0 DATA | @_UINT/CC/SCALbx34_ARA0 te=450-te-450 read args=0, E39                                                                           |
| 451 | 922 | R1 DATA | @_UINT/CC/SCALbx34_ARA0 te=451-te-451 read args=0, TCpr0.29_V_0                                                                  |
| 452 | 922 | R2 DATA |                                                                                                                                  |
| 452 | 922 | W0 DATA | EXEC ;@_UINT/CC/SCALbx36_crc_reg te=452-te-452 scalarw args=E40;@_UINT/CC/SCALbx36_byteno te=452-te-452 scalarw args=E41;TCpr0.\ |
|     |     |         | 35_V_0 te=452-te-452 scalarw args=E42 W/P:crc update hex:  reg...                                                                |
*-----+-----+---------+----------------------------------------------------------------------------------------------------------------------------------*

// res3: Thread=xpc10 state=X29:"29:xpc10:29"
*-----+-----+---------+---------------------------------------------------------------------------------------------------------------------------------------------------------*
| npc | eno | Phaser  | Work                                                                                                                                                    |
*-----+-----+---------+---------------------------------------------------------------------------------------------------------------------------------------------------------*
| 447 | -   | R0 CTRL |                                                                                                                                                         |
| 447 | 921 | R0 DATA | @_UINT/CC/SCALbx34_ARA0 te=447-te-447 read args=0, E37                                                                                                  |
| 448 | 921 | R1 DATA | @_UINT/CC/SCALbx34_ARA0 te=448-te-448 read args=0, TCpr0.35_V_0                                                                                         |
| 449 | 921 | R2 DATA |                                                                                                                                                         |
| 449 | 921 | W0 DATA | EXEC ;TSPcr2.16_V_1 te=449-te-449 scalarw args=C(1+TSPcr2.16_V_1);@_UINT/CC/SCALbx36_crc_reg te=449-te-449 scalarw args=E38 W/P:crc update hex:  reg... |
*-----+-----+---------+---------------------------------------------------------------------------------------------------------------------------------------------------------*

// res3: Thread=xpc10 state=X30:"30:xpc10:30"
*-----+-----+---------+-------------------------------------------------------------------*
| npc | eno | Phaser  | Work                                                              |
*-----+-----+---------+-------------------------------------------------------------------*
| 446 | -   | R0 CTRL |                                                                   |
| 446 | 919 | R0 DATA |                                                                   |
| 446 | 919 | W0 DATA | EXEC ;TSPte2.13_V_0 te=446-te-446 scalarw args=C(1+TSPte2.13_V_0) |
| 446 | 920 | R0 DATA |                                                                   |
| 446 | 920 | W0 DATA | EXEC                                                              |
*-----+-----+---------+-------------------------------------------------------------------*

// res3: Thread=xpc10 state=X31:"31:xpc10:31"
*-----+-----+---------+-----------------------------------------------------------------------------------------------*
| npc | eno | Phaser  | Work                                                                                          |
*-----+-----+---------+-----------------------------------------------------------------------------------------------*
| 442 | -   | R0 CTRL |                                                                                               |
| 442 | 918 | R0 DATA | iuMULTIPLIER14 te=442-te-442 *fixed-function-structural-alu* args=C64u(TSPte2.13_V_1), E2     |
| 443 | 918 | R1 DATA |                                                                                               |
| 444 | 918 | R2 DATA | @64_SS/CC/SCALbx54_ARB0 te=444-te-444 read args=0, E36                                        |
| 445 | 918 | R3 DATA |                                                                                               |
| 445 | 918 | W0 DATA | EXEC ;TSPte2.13_V_2 te=445-te-445 scalarw args=C(1+TSPte2.13_V_2) W/P:GSAI:hpr_writeln:$$A... |
*-----+-----+---------+-----------------------------------------------------------------------------------------------*

// res3: Thread=xpc10 state=X32:"32:xpc10:32"
*-----+-----+---------+-------------------------------------------------------------------------------------------------------------------------*
| npc | eno | Phaser  | Work                                                                                                                    |
*-----+-----+---------+-------------------------------------------------------------------------------------------------------------------------*
| 436 | -   | R0 CTRL | iuMULTIPLIER14 te=436-te-436 *fixed-function-structural-alu* args=C64u(TSPne2.10_V_0), E4;iuMULTIPLIER12 te=436-te-436\ |
|     |     |         |  *fixed-function-structural-alu* args=C64u(TSPne2.10_V_0), E3                                                           |
| 437 | -   | R1 CTRL |                                                                                                                         |
| 438 | -   | R2 CTRL | @64_SS/CC/SCALbx52_ARA0 te=438-te-438 read args=0, E31;@64_SS/CC/SCALbx58_ARD0 te=438-te-438 read args=0, E32           |
| 439 | -   | R3 CTRL |                                                                                                                         |
| 439 | 916 | R3 DATA |                                                                                                                         |
| 439 | 916 | W0 DATA | EXEC ;@64_SS/CC/SCALbx58_ARD0 te=439-te-439 write args=0, E29, E33;TSPne2.10_V_4 te=439-te-439 scalarw args=E34         |
| 440 | 916 | W1 DATA |                                                                                                                         |
| 439 | 917 | R3 DATA |                                                                                                                         |
| 439 | 917 | W0 DATA | EXEC ;@64_SS/CC/SCALbx58_ARD0 te=439-te-439 write args=0, E29, E35;TSPne2.10_V_4 te=439-te-439 scalarw args=E34         |
| 441 | 917 | W1 DATA |                                                                                                                         |
*-----+-----+---------+-------------------------------------------------------------------------------------------------------------------------*

// res3: Thread=xpc10 state=X33:"33:xpc10:33"
*-----+-----+---------+-------------------------------------------------------------------------------------------------------------------------*
| npc | eno | Phaser  | Work                                                                                                                    |
*-----+-----+---------+-------------------------------------------------------------------------------------------------------------------------*
| 430 | -   | R0 CTRL | iuMULTIPLIER14 te=430-te-430 *fixed-function-structural-alu* args=C64u(TSPne2.10_V_1), E1;iuMULTIPLIER12 te=430-te-430\ |
|     |     |         |  *fixed-function-structural-alu* args=C64u(TSPne2.10_V_1), E3                                                           |
| 431 | -   | R1 CTRL |                                                                                                                         |
| 432 | -   | R2 CTRL | @64_SS/CC/SCALbx52_ARA0 te=432-te-432 read args=0, E25;@64_SS/CC/SCALbx56_ARC0 te=432-te-432 read args=0, E26           |
| 433 | -   | R3 CTRL |                                                                                                                         |
| 433 | 914 | R3 DATA |                                                                                                                         |
| 433 | 914 | W0 DATA | EXEC ;@64_SS/CC/SCALbx56_ARC0 te=433-te-433 write args=0, E27, E28                                                      |
| 434 | 914 | W1 DATA |                                                                                                                         |
| 433 | 915 | R3 DATA |                                                                                                                         |
| 433 | 915 | W0 DATA | EXEC ;@64_SS/CC/SCALbx58_ARD0 te=433-te-433 write args=0, E29, E30                                                      |
| 435 | 915 | W1 DATA |                                                                                                                         |
*-----+-----+---------+-------------------------------------------------------------------------------------------------------------------------*

// res3: Thread=xpc10 state=X34:"34:xpc10:34"
*-----+-----+---------+-------------------------------------------------------------------------------------------------------------------------*
| npc | eno | Phaser  | Work                                                                                                                    |
*-----+-----+---------+-------------------------------------------------------------------------------------------------------------------------*
| 426 | -   | R0 CTRL | iuMULTIPLIER14 te=426-te-426 *fixed-function-structural-alu* args=C64u(TSPne2.10_V_0), E1;iuMULTIPLIER12 te=426-te-426\ |
|     |     |         |  *fixed-function-structural-alu* args=C64u(TSPne2.10_V_0), E4                                                           |
| 427 | -   | R1 CTRL |                                                                                                                         |
| 428 | -   | R2 CTRL | @64_SS/CC/SCALbx56_ARC0 te=428-te-428 read args=0, E21;@64_SS/CC/SCALbx58_ARD0 te=428-te-428 read args=0, E22           |
| 429 | -   | R3 CTRL |                                                                                                                         |
| 429 | 912 | R3 DATA |                                                                                                                         |
| 429 | 912 | W0 DATA | EXEC ;TSPne2.10_V_7 te=429-te-429 scalarw args=E23                                                                      |
| 429 | 913 | R3 DATA |                                                                                                                         |
| 429 | 913 | W0 DATA | EXEC ;TSPne2.10_V_7 te=429-te-429 scalarw args=E24                                                                      |
*-----+-----+---------+-------------------------------------------------------------------------------------------------------------------------*

// res3: Thread=xpc10 state=X35:"35:xpc10:35"
*-----+-----+---------+-------------------------------------------------------------------------------------------*
| npc | eno | Phaser  | Work                                                                                      |
*-----+-----+---------+-------------------------------------------------------------------------------------------*
| 422 | -   | R0 CTRL | iuMULTIPLIER14 te=422-te-422 *fixed-function-structural-alu* args=C64u(TSPne2.10_V_0), E2 |
| 423 | -   | R1 CTRL |                                                                                           |
| 424 | -   | R2 CTRL | @64_SS/CC/SCALbx54_ARB0 te=424-te-424 read args=0, E19                                    |
| 425 | -   | R3 CTRL |                                                                                           |
| 425 | 910 | R3 DATA |                                                                                           |
| 425 | 910 | W0 DATA | EXEC ;TSPne2.10_V_7 te=425-te-425 scalarw args=E20                                        |
| 425 | 911 | R3 DATA |                                                                                           |
| 425 | 911 | W0 DATA | EXEC                                                                                      |
*-----+-----+---------+-------------------------------------------------------------------------------------------*

// res3: Thread=xpc10 state=X36:"36:xpc10:36"
*-----+-----+---------+--------------------------------------------------------------------------------------------*
| npc | eno | Phaser  | Work                                                                                       |
*-----+-----+---------+--------------------------------------------------------------------------------------------*
| 416 | -   | R0 CTRL | iuMULTIPLIER14 te=416-te-416 *fixed-function-structural-alu* args=C64u(TSPne2.10_V_4), E16 |
| 417 | -   | R1 CTRL |                                                                                            |
| 418 | -   | R2 CTRL | @_SINT/CC/SCALbx16_ARA0 te=418-te-418 read args=0, E17                                     |
| 419 | -   | R3 CTRL |                                                                                            |
| 419 | 908 | R3 DATA |                                                                                            |
| 419 | 908 | W0 DATA | EXEC ;@64_SS/CC/SCALbx54_ARB0 te=419-te-419 write args=0, E13, C64(0)                      |
| 420 | 908 | W1 DATA |                                                                                            |
| 419 | 909 | R3 DATA |                                                                                            |
| 419 | 909 | W0 DATA | EXEC ;@64_SS/CC/SCALbx54_ARB0 te=419-te-419 write args=0, E13, E18                         |
| 421 | 909 | W1 DATA |                                                                                            |
*-----+-----+---------+--------------------------------------------------------------------------------------------*

// res3: Thread=xpc10 state=X37:"37:xpc10:37"
*-----+-----+---------+-------------------------------------------------------------------------------------------------------------------------*
| npc | eno | Phaser  | Work                                                                                                                    |
*-----+-----+---------+-------------------------------------------------------------------------------------------------------------------------*
| 411 | -   | R0 CTRL |                                                                                                                         |
| 411 | 907 | R0 DATA | iuMULTIPLIER14 te=411-te-411 *fixed-function-structural-alu* args=C64u(TSPne2.10_V_1), E2;iuMULTIPLIER12 te=411-te-411\ |
|     |     |         |  *fixed-function-structural-alu* args=C64u(TSPne2.10_V_1), E3                                                           |
| 412 | 907 | R1 DATA |                                                                                                                         |
| 413 | 907 | R2 DATA | @64_SS/CC/SCALbx54_ARB0 te=413-te-413 read args=0, E13                                                                  |
| 414 | 907 | R3 DATA |                                                                                                                         |
| 414 | 907 | W0 DATA | EXEC ;@64_SS/CC/SCALbx52_ARA0 te=414-te-414 write args=0, E14, E15;TSPne2.10_V_3 te=414-te-414 scalarw args=C(1+TSPne2\ |
|     |     |         | .10_V_3)                                                                                                                |
| 415 | 907 | W1 DATA |                                                                                                                         |
*-----+-----+---------+-------------------------------------------------------------------------------------------------------------------------*

// res3: Thread=xpc10 state=X38:"38:xpc10:38"
*-----+-----+---------+-----------------------------------------------------------------------------------------------------------------------------------*
| npc | eno | Phaser  | Work                                                                                                                              |
*-----+-----+---------+-----------------------------------------------------------------------------------------------------------------------------------*
| 409 | -   | R0 CTRL | @16_SS/CC/SCALbx10_ARA0 te=409-te-409 read args=0, TSPru0.12_V_1;@16_SS/CC/SCALbx12_ARB0 te=409-te-409 read args=0, TSPen0.17_V_0 |
| 410 | -   | R1 CTRL |                                                                                                                                   |
| 410 | 905 | R1 DATA |                                                                                                                                   |
| 410 | 905 | W0 DATA | EXEC ;TSPe0._SPILL_256 te=410-te-410 scalarw args=C(TSPen0.17_V_0)                                                                |
| 410 | 906 | R1 DATA |                                                                                                                                   |
| 410 | 906 | W0 DATA | EXEC ;TSPen0.17_V_0 te=410-te-410 scalarw args=C(1+TSPen0.17_V_0)                                                                 |
*-----+-----+---------+-----------------------------------------------------------------------------------------------------------------------------------*

// res3: Thread=xpc10 state=X39:"39:xpc10:39"
*-----+-----+---------+-----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------*
| npc | eno | Phaser  | Work                                                                                                                                                                                                                  |
*-----+-----+---------+-----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------*
| 407 | -   | R0 CTRL |                                                                                                                                                                                                                       |
| 407 | 904 | R0 DATA |                                                                                                                                                                                                                       |
| 407 | 904 | W0 DATA | EXEC ;@64_SS/CC/SCALbx52_ARA0 te=407-te-407 write args=0, E9, C64(-10);@64_SS/CC/SCALbx54_ARB0 te=407-te-407 write args=0, E10, C64(0);@64_SS/CC/SCALbx56_ARC0 te=407-te-407 write args=0, E11, C64(0);@64_SS/CC/SCA\ |
|     |     |         | Lbx58_ARD0 te=407-te-407 write args=0, E12, C64(0);TSPsw1.2_V_1 te=407-te-407 scalarw args=C(1+TSPsw1.2_V_1)                                                                                                          |
| 408 | 904 | W1 DATA |                                                                                                                                                                                                                       |
*-----+-----+---------+-----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------*

// res3: Thread=xpc10 state=X40:"40:xpc10:40"
*-----+-----+---------+----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------*
| npc | eno | Phaser  | Work                                                                                                                                                                                                                                                     |
*-----+-----+---------+----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------*
| 402 | -   | R0 CTRL |                                                                                                                                                                                                                                                          |
| 402 | 903 | R0 DATA | iuMULTIPLIER14 te=402-te-402 *fixed-function-structural-alu* args=C64u(TSPsw1.2_V_0), E1;iuMULTIPLIER12 te=402-te-402 *fixed-function-structural-alu* args=C64u(TSPsw1.2_V_0), E2;iuMULTIPLIER10 te=402-te-402 *fixed-function-structural-alu* args=C64\ |
|     |     |         | u(TSPsw1.2_V_0), E3                                                                                                                                                                                                                                      |
| 403 | 903 | R1 DATA | iuMULTIPLIER14 te=403-te-403 *fixed-function-structural-alu* args=C64u(TSPsw1.2_V_0), E4                                                                                                                                                                 |
| 404 | 903 | R2 DATA |                                                                                                                                                                                                                                                          |
| 405 | 903 | R3 DATA |                                                                                                                                                                                                                                                          |
| 405 | 903 | W0 DATA | EXEC ;TSPsw1.2_V_0 te=405-te-405 scalarw args=C(1+TSPsw1.2_V_0);d_monitor te=405-te-405 scalarw args=C64(TSPsw1.2_V_0);@64_SS/CC/SCALbx52_ARA0 te=405-te-405 write args=0, E5, C64(-10);@64_SS/CC/SCALbx54_ARB0 te=405-te-405 write args=0, E6, C64(0);\ |
|     |     |         | @64_SS/CC/SCALbx56_ARC0 te=405-te-405 write args=0, E7, C64(0);@64_SS/CC/SCALbx58_ARD0 te=405-te-405 write args=0, E8, C64(0)                                                                                                                            |
| 406 | 903 | W1 DATA |                                                                                                                                                                                                                                                          |
*-----+-----+---------+----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------*

// res3: Thread=xpc10 state=X41:"41:xpc10:41"
*-----+-----+---------+--------------------------------------------------------*
| npc | eno | Phaser  | Work                                                   |
*-----+-----+---------+--------------------------------------------------------*
| 401 | -   | R0 CTRL |                                                        |
| 401 | 901 | R0 DATA |                                                        |
| 401 | 901 | W0 DATA | EXEC ;TSPe1._SPILL_256 te=401-te-401 scalarw args=C(0) |
| 401 | 902 | R0 DATA |                                                        |
| 401 | 902 | W0 DATA | EXEC                                                   |
*-----+-----+---------+--------------------------------------------------------*

// res3: Thread=xpc10 state=X0:"0:xpc10:start0"
*-----+-----+-----------+--------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------*
| npc | eno | Phaser    | Work                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   |
*-----+-----+-----------+--------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------*
| 0   | -   | R0 CTRL   |                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        |
| 0   | 900 | R0 DATA   |                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        |
| 0   | 900 | W0 DATA   | EXEC ;TSPen1.8_V_0 te=0-te-0 scalarw args=C(0);TSPin0.6_V_0 te=0-te-0 scalarw args=C(0);phase te=0-te-0 scalarw args=Cu(2);@_SINT/CC/SCALbx40_d2dim0 te=0-te-0 scalarw args=C(78);@_SINT/CC/SCALbx42_d2dim0 te=0-te-0 scalarw args=C(78);@_SINT/CC/SCALbx44_d2dim0 te=0-te-0 scalarw args=C(78);@_SINT/CC/SCALbx46_d2dim0 te=0-te-0 scalarw args=C(78);@_SINT/CC/SCALbx32_d2dim0 te=0-te-0 scalarw args=C64(20);@_UINT/CC/SCALbx34_ARA0 te=0-te-0 write args=0, 255, Cu(-1309196108);@_SINT/CC/SCALbx\ |
|     |     |           | 16_ARA0 te=0-te-0 write args=0, 399, C(10);@16_SS/CC/SCALbx10_ARA0 te=0-te-0 write args=0, 74, C16(108);@16_SS/CC/SCALbx14_ARC0 te=0-te-0 write args=0, 76, C16(110);@16_SS/CC/SCALbx12_ARB0 te=0-te-0 write args=0, 19, C16(121) W/P:waypoint %u %u                                                                                                                                                                                                                                                   |
| 1   | 900 | W1 DATA   | @_UINT/CC/SCALbx34_ARA0 te=1-te-1 write args=0, 254, Cu(-1254728445);@_SINT/CC/SCALbx16_ARA0 te=1-te-1 write args=0, 398, C(0);@16_SS/CC/SCALbx10_ARA0 te=1-te-1 write args=0, 73, C16(112);@16_SS/CC/SCALbx14_ARC0 te=1-te-1 write args=0, 75, C16(101);@16_SS/CC/SCALbx12_ARB0 te=1-te-1 write args=0, 18, C16(119)                                                                                                                                                                                  |
| 2   | 900 | W2 DATA   | @_UINT/CC/SCALbx34_ARA0 te=2-te-2 write args=0, 253, Cu(-1200260134);@_SINT/CC/SCALbx16_ARA0 te=2-te-2 write args=0, 397, C(-2);@16_SS/CC/SCALbx10_ARA0 te=2-te-2 write args=0, 72, C16(105);@16_SS/CC/SCALbx14_ARC0 te=2-te-2 write args=0, 74, C16(113);@16_SS/CC/SCALbx12_ARB0 te=2-te-2 write args=0, 17, C16(118)                                                                                                                                                                                 |
| 3   | 900 | W3 DATA   | @_UINT/CC/SCALbx34_ARA0 te=3-te-3 write args=0, 252, Cu(-1129027987);@_SINT/CC/SCALbx16_ARA0 te=3-te-3 write args=0, 396, C(-3);@16_SS/CC/SCALbx10_ARA0 te=3-te-3 write args=0, 71, C16(116);@16_SS/CC/SCALbx14_ARC0 te=3-te-3 write args=0, 73, C16(114);@16_SS/CC/SCALbx12_ARB0 te=3-te-3 write args=0, 16, C16(116)                                                                                                                                                                                 |
| 4   | 900 | W4 DATA   | @_UINT/CC/SCALbx34_ARA0 te=4-te-4 write args=0, 251, Cu(-1561119128);@_SINT/CC/SCALbx16_ARA0 te=4-te-4 write args=0, 395, C(-3);@16_SS/CC/SCALbx10_ARA0 te=4-te-4 write args=0, 70, C16(101);@16_SS/CC/SCALbx14_ARC0 te=4-te-4 write args=0, 72, C16(118);@16_SS/CC/SCALbx12_ARB0 te=4-te-4 write args=0, 15, C16(115)                                                                                                                                                                                 |
| 5   | 900 | W5 DATA   | @_UINT/CC/SCALbx34_ARA0 te=5-te-5 write args=0, 250, Cu(-1506661409);@_SINT/CC/SCALbx16_ARA0 te=5-te-5 write args=0, 394, C(-4);@16_SS/CC/SCALbx10_ARA0 te=5-te-5 write args=0, 69, C16(121);@16_SS/CC/SCALbx14_ARC0 te=5-te-5 write args=0, 71, C16(101);@16_SS/CC/SCALbx12_ARB0 te=5-te-5 write args=0, 14, C16(114)                                                                                                                                                                                 |
| 6   | 900 | W6 DATA   | @_UINT/CC/SCALbx34_ARA0 te=6-te-6 write args=0, 249, Cu(-1418654458);@_SINT/CC/SCALbx16_ARA0 te=6-te-6 write args=0, 393, C(-4);@16_SS/CC/SCALbx10_ARA0 te=6-te-6 write args=0, 68, C16(103);@16_SS/CC/SCALbx14_ARC0 te=6-te-6 write args=0, 70, C16(107);@16_SS/CC/SCALbx12_ARB0 te=6-te-6 write args=0, 13, C16(113)                                                                                                                                                                                 |
| 7   | 900 | W7 DATA   | @_UINT/CC/SCALbx34_ARA0 te=7-te-7 write args=0, 248, Cu(-1347415887);@_SINT/CC/SCALbx16_ARA0 te=7-te-7 write args=0, 392, C(-5);@16_SS/CC/SCALbx10_ARA0 te=7-te-7 write args=0, 67, C16(113);@16_SS/CC/SCALbx14_ARC0 te=7-te-7 write args=0, 69, C16(97);@16_SS/CC/SCALbx12_ARB0 te=7-te-7 write args=0, 12, C16(112)                                                                                                                                                                                  |
| 8   | 900 | W8 DATA   | @_UINT/CC/SCALbx34_ARA0 te=8-te-8 write args=0, 247, Cu(-1744851700);@_SINT/CC/SCALbx16_ARA0 te=8-te-8 write args=0, 391, C(-2);@16_SS/CC/SCALbx10_ARA0 te=8-te-8 write args=0, 66, C16(105);@16_SS/CC/SCALbx14_ARC0 te=8-te-8 write args=0, 68, C16(101);@16_SS/CC/SCALbx12_ARB0 te=8-te-8 write args=0, 11, C16(110)                                                                                                                                                                                 |
| 9   | 900 | W9 DATA   | @_UINT/CC/SCALbx34_ARA0 te=9-te-9 write args=0, 246, Cu(-1824608069);@_SINT/CC/SCALbx16_ARA0 te=9-te-9 write args=0, 390, C(-2);@16_SS/CC/SCALbx10_ARA0 te=9-te-9 write args=0, 65, C16(114);@16_SS/CC/SCALbx14_ARC0 te=9-te-9 write args=0, 67, C16(101);@16_SS/CC/SCALbx12_ARB0 te=9-te-9 write args=0, 10, C16(109)                                                                                                                                                                                 |
| 10  | 900 | W10 DATA  | @_UINT/CC/SCALbx34_ARA0 te=10-te-10 write args=0, 245, Cu(-1635936670);@_SINT/CC/SCALbx16_ARA0 te=10-te-10 write args=0, 389, C(-1);@16_SS/CC/SCALbx10_ARA0 te=10-te-10 write args=0, 64, C16(97);@16_SS/CC/SCALbx14_ARC0 te=10-te-10 write args=0, 66, C16(108);@16_SS/CC/SCALbx12_ARB0 te=10-te-10 write args=0, 9, C16(108)                                                                                                                                                                         |
| 11  | 900 | W11 DATA  | @_UINT/CC/SCALbx34_ARA0 te=11-te-11 write args=0, 244, Cu(-1698919467);@_SINT/CC/SCALbx16_ARA0 te=11-te-11 write args=0, 388, C(-4);@16_SS/CC/SCALbx10_ARA0 te=11-te-11 write args=0, 63, C16(118);@16_SS/CC/SCALbx14_ARC0 te=11-te-11 write args=0, 65, C16(97);@16_SS/CC/SCALbx12_ARB0 te=11-te-11 write args=0, 8, C16(107)                                                                                                                                                                         |
| 12  | 900 | W12 DATA  | @_UINT/CC/SCALbx34_ARA0 te=12-te-12 write args=0, 243, Cu(-2063868976);@_SINT/CC/SCALbx16_ARA0 te=12-te-12 write args=0, 387, C(-1);@16_SS/CC/SCALbx10_ARA0 te=12-te-12 write args=0, 62, C16(101);@16_SS/CC/SCALbx14_ARC0 te=12-te-12 write args=0, 64, C16(101);@16_SS/CC/SCALbx12_ARB0 te=12-te-12 write args=0, 7, C16(105)                                                                                                                                                                        |
| 13  | 900 | W13 DATA  | @_UINT/CC/SCALbx34_ARA0 te=13-te-13 write args=0, 242, Cu(-2143631769);@_SINT/CC/SCALbx16_ARA0 te=13-te-13 write args=0, 386, C(0);@16_SS/CC/SCALbx10_ARA0 te=13-te-13 write args=0, 61, C16(101);@16_SS/CC/SCALbx14_ARC0 te=13-te-13 write args=0, 63, C16(113);@16_SS/CC/SCALbx12_ARB0 te=13-te-13 write args=0, 6, C16(104)                                                                                                                                                                         |
| 14  | 900 | W14 DATA  | @_UINT/CC/SCALbx34_ARA0 te=14-te-14 write args=0, 241, Cu(-1921392450);@_SINT/CC/SCALbx16_ARA0 te=14-te-14 write args=0, 385, C(-5);@16_SS/CC/SCALbx10_ARA0 te=14-te-14 write args=0, 60, C16(118);@16_SS/CC/SCALbx14_ARC0 te=14-te-14 write args=0, 62, C16(115);@16_SS/CC/SCALbx12_ARB0 te=14-te-14 write args=0, 5, C16(103)                                                                                                                                                                        |
| 15  | 900 | W15 DATA  | @_UINT/CC/SCALbx34_ARA0 te=15-te-15 write args=0, 240, Cu(-1984365303);@_SINT/CC/SCALbx16_ARA0 te=15-te-15 write args=0, 384, C(7);@16_SS/CC/SCALbx10_ARA0 te=15-te-15 write args=0, 59, C16(108);@16_SS/CC/SCALbx14_ARC0 te=15-te-15 write args=0, 61, C16(103);@16_SS/CC/SCALbx12_ARB0 te=15-te-15 write args=0, 4, C16(102)                                                                                                                                                                         |
| 16  | 900 | W16 DATA  | @_UINT/CC/SCALbx34_ARA0 te=16-te-16 write args=0, 239, Cu(-35218492);@_SINT/CC/SCALbx16_ARA0 te=16-te-16 write args=0, 383, C(-4);@16_SS/CC/SCALbx10_ARA0 te=16-te-16 write args=0, 58, C16(100);@16_SS/CC/SCALbx14_ARC0 te=16-te-16 write args=0, 60, C16(119);@16_SS/CC/SCALbx12_ARB0 te=16-te-16 write args=0, 3, C16(101)                                                                                                                                                                          |
| 17  | 900 | W17 DATA  | @_UINT/CC/SCALbx34_ARA0 te=17-te-17 write args=0, 238, Cu(-114850189);@_SINT/CC/SCALbx16_ARA0 te=17-te-17 write args=0, 382, C(-4);@16_SS/CC/SCALbx10_ARA0 te=17-te-17 write args=0, 57, C16(101);@16_SS/CC/SCALbx14_ARC0 te=17-te-17 write args=0, 59, C16(118);@16_SS/CC/SCALbx12_ARB0 te=17-te-17 write args=0, 2, C16(100)                                                                                                                                                                         |
| 18  | 900 | W18 DATA  | @_UINT/CC/SCALbx34_ARA0 te=18-te-18 write args=0, 237, Cu(-194731862);@_SINT/CC/SCALbx16_ARA0 te=18-te-18 write args=0, 381, C(0);@16_SS/CC/SCALbx10_ARA0 te=18-te-18 write args=0, 56, C16(101);@16_SS/CC/SCALbx14_ARC0 te=18-te-18 write args=0, 58, C16(101);@16_SS/CC/SCALbx12_ARB0 te=18-te-18 write args=0, 1, C16(99)                                                                                                                                                                           |
| 19  | 900 | W19 DATA  | @_UINT/CC/SCALbx34_ARA0 te=19-te-19 write args=0, 236, Cu(-257573603);@_SINT/CC/SCALbx16_ARA0 te=19-te-19 write args=0, 380, C(-3);@16_SS/CC/SCALbx10_ARA0 te=19-te-19 write args=0, 55, C16(108);@16_SS/CC/SCALbx14_ARC0 te=19-te-19 write args=0, 57, C16(108);@16_SS/CC/SCALbx12_ARB0 te=19-te-19 write args=0, 0, C16(97)                                                                                                                                                                          |
| 20  | 900 | W20 DATA  | @_UINT/CC/SCALbx34_ARA0 te=20-te-20 write args=0, 235, Cu(-287118056);@_SINT/CC/SCALbx16_ARA0 te=20-te-20 write args=0, 379, C(0);@16_SS/CC/SCALbx10_ARA0 te=20-te-20 write args=0, 54, C16(114);@16_SS/CC/SCALbx14_ARC0 te=20-te-20 write args=0, 56, C16(115)                                                                                                                                                                                                                                        |
| 21  | 900 | W21 DATA  | @_UINT/CC/SCALbx34_ARA0 te=21-te-21 write args=0, 234, Cu(-366743377);@_SINT/CC/SCALbx16_ARA0 te=21-te-21 write args=0, 378, C(17);@16_SS/CC/SCALbx10_ARA0 te=21-te-21 write args=0, 53, C16(108);@16_SS/CC/SCALbx14_ARC0 te=21-te-21 write args=0, 55, C16(114)                                                                                                                                                                                                                                       |
| 22  | 900 | W22 DATA  | @_UINT/CC/SCALbx34_ARA0 te=22-te-22 write args=0, 233, Cu(-413084042);@_SINT/CC/SCALbx16_ARA0 te=22-te-22 write args=0, 377, C(-6);@16_SS/CC/SCALbx10_ARA0 te=22-te-22 write args=0, 52, C16(100);@16_SS/CC/SCALbx14_ARC0 te=22-te-22 write args=0, 54, C16(107)                                                                                                                                                                                                                                       |
| 23  | 900 | W23 DATA  | @_UINT/CC/SCALbx34_ARA0 te=23-te-23 write args=0, 232, Cu(-475935807);@_SINT/CC/SCALbx16_ARA0 te=23-te-23 write args=0, 376, C(-5);@16_SS/CC/SCALbx10_ARA0 te=23-te-23 write args=0, 51, C16(108);@16_SS/CC/SCALbx14_ARC0 te=23-te-23 write args=0, 53, C16(118)                                                                                                                                                                                                                                       |
| 24  | 900 | W24 DATA  | @_UINT/CC/SCALbx34_ARA0 te=24-te-24 write args=0, 231, Cu(-605129092);@_SINT/CC/SCALbx16_ARA0 te=24-te-24 write args=0, 375, C(-2);@16_SS/CC/SCALbx10_ARA0 te=24-te-24 write args=0, 50, C16(114);@16_SS/CC/SCALbx14_ARC0 te=24-te-24 write args=0, 52, C16(105)                                                                                                                                                                                                                                       |
| 25  | 900 | W25 DATA  | @_UINT/CC/SCALbx34_ARA0 te=25-te-25 write args=0, 230, Cu(-550540341);@_SINT/CC/SCALbx16_ARA0 te=25-te-25 write args=0, 374, C(2);@16_SS/CC/SCALbx10_ARA0 te=25-te-25 write args=0, 49, C16(104);@16_SS/CC/SCALbx14_ARC0 te=25-te-25 write args=0, 51, C16(113)                                                                                                                                                                                                                                        |
| 26  | 900 | W26 DATA  | @_UINT/CC/SCALbx34_ARA0 te=26-te-26 write args=0, 229, Cu(-764654318);@_SINT/CC/SCALbx16_ARA0 te=26-te-26 write args=0, 373, C(-5);@16_SS/CC/SCALbx10_ARA0 te=26-te-26 write args=0, 48, C16(115);@16_SS/CC/SCALbx14_ARC0 te=26-te-26 write args=0, 50, C16(108)                                                                                                                                                                                                                                       |
| 27  | 900 | W27 DATA  | @_UINT/CC/SCALbx34_ARA0 te=27-te-27 write args=0, 228, Cu(-693284699);@_SINT/CC/SCALbx16_ARA0 te=27-te-27 write args=0, 372, C(-6);@16_SS/CC/SCALbx10_ARA0 te=27-te-27 write args=0, 47, C16(112);@16_SS/CC/SCALbx14_ARC0 te=27-te-27 write args=0, 49, C16(107)                                                                                                                                                                                                                                       |
| 28  | 900 | W28 DATA  | @_UINT/CC/SCALbx34_ARA0 te=28-te-28 write args=0, 227, Cu(-924188512);@_SINT/CC/SCALbx16_ARA0 te=28-te-28 write args=0, 371, C(-4);@16_SS/CC/SCALbx10_ARA0 te=28-te-28 write args=0, 46, C16(112);@16_SS/CC/SCALbx14_ARC0 te=28-te-28 write args=0, 48, C16(108)                                                                                                                                                                                                                                       |
| 29  | 900 | W29 DATA  | @_UINT/CC/SCALbx34_ARA0 te=29-te-29 write args=0, 226, Cu(-869589737);@_SINT/CC/SCALbx16_ARA0 te=29-te-29 write args=0, 370, C(-4);@16_SS/CC/SCALbx10_ARA0 te=29-te-29 write args=0, 45, C16(116);@16_SS/CC/SCALbx14_ARC0 te=29-te-29 write args=0, 47, C16(121)                                                                                                                                                                                                                                       |
| 30  | 900 | W30 DATA  | @_UINT/CC/SCALbx34_ARA0 te=30-te-30 write args=0, 225, Cu(-1050133554);@_SINT/CC/SCALbx16_ARA0 te=30-te-30 write args=0, 369, C(-2);@16_SS/CC/SCALbx10_ARA0 te=30-te-30 write args=0, 44, C16(118);@16_SS/CC/SCALbx14_ARC0 te=30-te-30 write args=0, 46, C16(108)                                                                                                                                                                                                                                      |
| 31  | 900 | W31 DATA  | @_UINT/CC/SCALbx34_ARA0 te=31-te-31 write args=0, 224, Cu(-978770311);@_SINT/CC/SCALbx16_ARA0 te=31-te-31 write args=0, 368, C(-3);@16_SS/CC/SCALbx10_ARA0 te=31-te-31 write args=0, 43, C16(114);@16_SS/CC/SCALbx14_ARC0 te=31-te-31 write args=0, 45, C16(107)                                                                                                                                                                                                                                       |
| 32  | 900 | W32 DATA  | @_UINT/CC/SCALbx34_ARA0 te=32-te-32 write args=0, 223, Cu(701822548);@_SINT/CC/SCALbx16_ARA0 te=32-te-32 write args=0, 367, C(-5);@16_SS/CC/SCALbx10_ARA0 te=32-te-32 write args=0, 42, C16(121);@16_SS/CC/SCALbx14_ARC0 te=32-te-32 write args=0, 44, C16(109)                                                                                                                                                                                                                                        |
| 33  | 900 | W33 DATA  | @_UINT/CC/SCALbx34_ARA0 te=33-te-33 write args=0, 222, Cu(756411363);@_SINT/CC/SCALbx16_ARA0 te=33-te-33 write args=0, 366, C(-3);@16_SS/CC/SCALbx10_ARA0 te=33-te-33 write args=0, 41, C16(116);@16_SS/CC/SCALbx14_ARC0 te=33-te-33 write args=0, 43, C16(100)                                                                                                                                                                                                                                        |
| 34  | 900 | W34 DATA  | @_UINT/CC/SCALbx34_ARA0 te=34-te-34 write args=0, 221, Cu(542559546);@_SINT/CC/SCALbx16_ARA0 te=34-te-34 write args=0, 365, C(-7);@16_SS/CC/SCALbx10_ARA0 te=34-te-34 write args=0, 40, C16(112);@16_SS/CC/SCALbx14_ARC0 te=34-te-34 write args=0, 42, C16(103)                                                                                                                                                                                                                                        |
| 35  | 900 | W35 DATA  | @_UINT/CC/SCALbx34_ARA0 te=35-te-35 write args=0, 220, Cu(613929101);@_SINT/CC/SCALbx16_ARA0 te=35-te-35 write args=0, 364, C(0);@16_SS/CC/SCALbx10_ARA0 te=35-te-35 write args=0, 39, C16(103);@16_SS/CC/SCALbx14_ARC0 te=35-te-35 write args=0, 41, C16(119)                                                                                                                                                                                                                                         |
| 36  | 900 | W36 DATA  | @_UINT/CC/SCALbx34_ARA0 te=36-te-36 write args=0, 219, Cu(986742920);@_SINT/CC/SCALbx16_ARA0 te=36-te-36 write args=0, 363, C(-7);@16_SS/CC/SCALbx10_ARA0 te=36-te-36 write args=0, 38, C16(101);@16_SS/CC/SCALbx14_ARC0 te=36-te-36 write args=0, 40, C16(113)                                                                                                                                                                                                                                        |
| 37  | 900 | W37 DATA  | @_UINT/CC/SCALbx34_ARA0 te=37-te-37 write args=0, 218, Cu(1041341759);@_SINT/CC/SCALbx16_ARA0 te=37-te-37 write args=0, 362, C(-7);@16_SS/CC/SCALbx10_ARA0 te=37-te-37 write args=0, 37, C16(103);@16_SS/CC/SCALbx14_ARC0 te=37-te-37 write args=0, 39, C16(115)                                                                                                                                                                                                                                       |
| 38  | 900 | W38 DATA  | @_UINT/CC/SCALbx34_ARA0 te=38-te-38 write args=0, 217, Cu(861060070);@_SINT/CC/SCALbx16_ARA0 te=38-te-38 write args=0, 361, C(-8);@16_SS/CC/SCALbx10_ARA0 te=38-te-38 write args=0, 36, C16(101);@16_SS/CC/SCALbx14_ARC0 te=38-te-38 write args=0, 38, C16(104)                                                                                                                                                                                                                                        |
| 39  | 900 | W39 DATA  | @_UINT/CC/SCALbx34_ARA0 te=39-te-39 write args=0, 216, Cu(932423249);@_SINT/CC/SCALbx16_ARA0 te=39-te-39 write args=0, 360, C(-6);@16_SS/CC/SCALbx10_ARA0 te=39-te-39 write args=0, 35, C16(118);@16_SS/CC/SCALbx14_ARC0 te=39-te-39 write args=0, 37, C16(104)                                                                                                                                                                                                                                        |
| 40  | 900 | W40 DATA  | @_UINT/CC/SCALbx34_ARA0 te=40-te-40 write args=0, 215, Cu(266083308);@_SINT/CC/SCALbx16_ARA0 te=40-te-40 write args=0, 359, C(-2);@16_SS/CC/SCALbx10_ARA0 te=40-te-40 write args=0, 34, C16(114);@16_SS/CC/SCALbx14_ARC0 te=40-te-40 write args=0, 36, C16(112)                                                                                                                                                                                                                                        |
| 41  | 900 | W41 DATA  | @_UINT/CC/SCALbx34_ARA0 te=41-te-41 write args=0, 214, Cu(186451547);@_SINT/CC/SCALbx16_ARA0 te=41-te-41 write args=0, 358, C(-6);@16_SS/CC/SCALbx10_ARA0 te=41-te-41 write args=0, 33, C16(99);@16_SS/CC/SCALbx14_ARC0 te=41-te-41 write args=0, 35, C16(110)                                                                                                                                                                                                                                         |
| 42  | 900 | W42 DATA  | @_UINT/CC/SCALbx34_ARA0 te=42-te-42 write args=0, 213, Cu(106832002);@_SINT/CC/SCALbx16_ARA0 te=42-te-42 write args=0, 357, C(4);@16_SS/CC/SCALbx10_ARA0 te=42-te-42 write args=0, 32, C16(103);@16_SS/CC/SCALbx14_ARC0 te=42-te-42 write args=0, 34, C16(107)                                                                                                                                                                                                                                         |
| 43  | 900 | W43 DATA  | @_UINT/CC/SCALbx34_ARA0 te=43-te-43 write args=0, 212, Cu(43990325);@_SINT/CC/SCALbx16_ARA0 te=43-te-43 write args=0, 356, C(0);@16_SS/CC/SCALbx10_ARA0 te=43-te-43 write args=0, 31, C16(108);@16_SS/CC/SCALbx14_ARC0 te=43-te-43 write args=0, 33, C16(107)                                                                                                                                                                                                                                          |
| 44  | 900 | W44 DATA  | @_UINT/CC/SCALbx34_ARA0 te=44-te-44 write args=0, 211, Cu(483945776);@_SINT/CC/SCALbx16_ARA0 te=44-te-44 write args=0, 355, C(-1);@16_SS/CC/SCALbx10_ARA0 te=44-te-44 write args=0, 30, C16(114);@16_SS/CC/SCALbx14_ARC0 te=44-te-44 write args=0, 32, C16(118)                                                                                                                                                                                                                                        |
| 45  | 900 | W45 DATA  | @_UINT/CC/SCALbx34_ARA0 te=45-te-45 write args=0, 210, Cu(404320391);@_SINT/CC/SCALbx16_ARA0 te=45-te-45 write args=0, 354, C(-2);@16_SS/CC/SCALbx10_ARA0 te=45-te-45 write args=0, 29, C16(107);@16_SS/CC/SCALbx14_ARC0 te=45-te-45 write args=0, 31, C16(105)                                                                                                                                                                                                                                        |
| 46  | 900 | W46 DATA  | @_UINT/CC/SCALbx34_ARA0 te=46-te-46 write args=0, 209, Cu(358241886);@_SINT/CC/SCALbx16_ARA0 te=46-te-46 write args=0, 353, C(-2);@16_SS/CC/SCALbx10_ARA0 te=46-te-46 write args=0, 28, C16(108);@16_SS/CC/SCALbx14_ARC0 te=46-te-46 write args=0, 30, C16(102)                                                                                                                                                                                                                                        |
| 47  | 900 | W47 DATA  | @_UINT/CC/SCALbx34_ARA0 te=47-te-47 write args=0, 208, Cu(295390185);@_SINT/CC/SCALbx16_ARA0 te=47-te-47 write args=0, 352, C(-1);@16_SS/CC/SCALbx10_ARA0 te=47-te-47 write args=0, 27, C16(105);@16_SS/CC/SCALbx14_ARC0 te=47-te-47 write args=0, 29, C16(107)                                                                                                                                                                                                                                        |
| 48  | 900 | W48 DATA  | @_UINT/CC/SCALbx34_ARA0 te=48-te-48 write args=0, 207, Cu(1707420964);@_SINT/CC/SCALbx16_ARA0 te=48-te-48 write args=0, 351, C(-2);@16_SS/CC/SCALbx10_ARA0 te=48-te-48 write args=0, 26, C16(97);@16_SS/CC/SCALbx14_ARC0 te=48-te-48 write args=0, 28, C16(108)                                                                                                                                                                                                                                        |
| 49  | 900 | W49 DATA  | @_UINT/CC/SCALbx34_ARA0 te=49-te-49 write args=0, 206, Cu(1627664531);@_SINT/CC/SCALbx16_ARA0 te=49-te-49 write args=0, 350, C(2);@16_SS/CC/SCALbx10_ARA0 te=49-te-49 write args=0, 25, C16(105);@16_SS/CC/SCALbx14_ARC0 te=49-te-49 write args=0, 27, C16(112)                                                                                                                                                                                                                                        |
| 50  | 900 | W50 DATA  | @_UINT/CC/SCALbx34_ARA0 te=50-te-50 write args=0, 205, Cu(1816598090);@_SINT/CC/SCALbx16_ARA0 te=50-te-50 write args=0, 349, C(2);@16_SS/CC/SCALbx10_ARA0 te=50-te-50 write args=0, 24, C16(113);@16_SS/CC/SCALbx14_ARC0 te=50-te-50 write args=0, 26, C16(112)                                                                                                                                                                                                                                        |
| 51  | 900 | W51 DATA  | @_UINT/CC/SCALbx34_ARA0 te=51-te-51 write args=0, 204, Cu(1753615357);@_SINT/CC/SCALbx16_ARA0 te=51-te-51 write args=0, 348, C(-2);@16_SS/CC/SCALbx10_ARA0 te=51-te-51 write args=0, 23, C16(101);@16_SS/CC/SCALbx14_ARC0 te=51-te-51 write args=0, 25, C16(101)                                                                                                                                                                                                                                       |
| 52  | 900 | W52 DATA  | @_UINT/CC/SCALbx34_ARA0 te=52-te-52 write args=0, 203, Cu(1992383480);@_SINT/CC/SCALbx16_ARA0 te=52-te-52 write args=0, 347, C(4);@16_SS/CC/SCALbx10_ARA0 te=52-te-52 write args=0, 22, C16(97);@16_SS/CC/SCALbx14_ARC0 te=52-te-52 write args=0, 24, C16(114)                                                                                                                                                                                                                                         |
| 53  | 900 | W53 DATA  | @_UINT/CC/SCALbx34_ARA0 te=53-te-53 write args=0, 202, Cu(1912620623);@_SINT/CC/SCALbx16_ARA0 te=53-te-53 write args=0, 346, C(-2);@16_SS/CC/SCALbx10_ARA0 te=53-te-53 write args=0, 21, C16(101);@16_SS/CC/SCALbx14_ARC0 te=53-te-53 write args=0, 23, C16(107)                                                                                                                                                                                                                                       |
| 54  | 900 | W54 DATA  | @_UINT/CC/SCALbx34_ARA0 te=54-te-54 write args=0, 201, Cu(2135122070);@_SINT/CC/SCALbx16_ARA0 te=54-te-54 write args=0, 345, C(-1);@16_SS/CC/SCALbx10_ARA0 te=54-te-54 write args=0, 20, C16(112);@16_SS/CC/SCALbx14_ARC0 te=54-te-54 write args=0, 22, C16(101)                                                                                                                                                                                                                                       |
| 55  | 900 | W55 DATA  | @_UINT/CC/SCALbx34_ARA0 te=55-te-55 write args=0, 200, Cu(2072149281);@_SINT/CC/SCALbx16_ARA0 te=55-te-55 write args=0, 344, C(-1);@16_SS/CC/SCALbx10_ARA0 te=55-te-55 write args=0, 19, C16(121);@16_SS/CC/SCALbx14_ARC0 te=55-te-55 write args=0, 21, C16(108)                                                                                                                                                                                                                                       |
| 56  | 900 | W56 DATA  | @_UINT/CC/SCALbx34_ARA0 te=56-te-56 write args=0, 199, Cu(1137557660);@_SINT/CC/SCALbx16_ARA0 te=56-te-56 write args=0, 343, C(-2);@16_SS/CC/SCALbx10_ARA0 te=56-te-56 write args=0, 18, C16(115);@16_SS/CC/SCALbx14_ARC0 te=56-te-56 write args=0, 20, C16(100)                                                                                                                                                                                                                                       |
| 57  | 900 | W57 DATA  | @_UINT/CC/SCALbx34_ARA0 te=57-te-57 write args=0, 198, Cu(1192025387);@_SINT/CC/SCALbx16_ARA0 te=57-te-57 write args=0, 342, C(-2);@16_SS/CC/SCALbx10_ARA0 te=57-te-57 write args=0, 17, C16(116);@16_SS/CC/SCALbx14_ARC0 te=57-te-57 write args=0, 19, C16(99)                                                                                                                                                                                                                                        |
| 58  | 900 | W58 DATA  | @_UINT/CC/SCALbx34_ARA0 te=58-te-58 write args=0, 197, Cu(1246755826);@_SINT/CC/SCALbx16_ARA0 te=58-te-58 write args=0, 341, C(-2);@16_SS/CC/SCALbx10_ARA0 te=58-te-58 write args=0, 16, C16(103);@16_SS/CC/SCALbx14_ARC0 te=58-te-58 write args=0, 18, C16(100)                                                                                                                                                                                                                                       |
| 59  | 900 | W59 DATA  | @_UINT/CC/SCALbx34_ARA0 te=59-te-59 write args=0, 196, Cu(1317987909);@_SINT/CC/SCALbx16_ARA0 te=59-te-59 write args=0, 340, C(0);@16_SS/CC/SCALbx10_ARA0 te=59-te-59 write args=0, 15, C16(108);@16_SS/CC/SCALbx14_ARC0 te=59-te-59 write args=0, 17, C16(107)                                                                                                                                                                                                                                        |
| 60  | 900 | W60 DATA  | @_UINT/CC/SCALbx34_ARA0 te=60-te-60 write args=0, 195, Cu(1355396672);@_SINT/CC/SCALbx16_ARA0 te=60-te-60 write args=0, 339, C(-3);@16_SS/CC/SCALbx10_ARA0 te=60-te-60 write args=0, 14, C16(108);@16_SS/CC/SCALbx14_ARC0 te=60-te-60 write args=0, 16, C16(108)                                                                                                                                                                                                                                       |
| 61  | 900 | W61 DATA  | @_UINT/CC/SCALbx34_ARA0 te=61-te-61 write args=0, 194, Cu(1409854455);@_SINT/CC/SCALbx16_ARA0 te=61-te-61 write args=0, 338, C(-5);@16_SS/CC/SCALbx10_ARA0 te=61-te-61 write args=0, 13, C16(114);@16_SS/CC/SCALbx14_ARC0 te=61-te-61 write args=0, 15, C16(108)                                                                                                                                                                                                                                       |
| 62  | 900 | W62 DATA  | @_UINT/CC/SCALbx34_ARA0 te=62-te-62 write args=0, 193, Cu(1498123566);@_SINT/CC/SCALbx16_ARA0 te=62-te-62 write args=0, 337, C(0);@16_SS/CC/SCALbx10_ARA0 te=62-te-62 write args=0, 12, C16(110);@16_SS/CC/SCALbx14_ARC0 te=62-te-62 write args=0, 14, C16(121)                                                                                                                                                                                                                                        |
| 63  | 900 | W63 DATA  | @_UINT/CC/SCALbx34_ARA0 te=63-te-63 write args=0, 192, Cu(1569362073);@_SINT/CC/SCALbx16_ARA0 te=63-te-63 write args=0, 336, C(3);@16_SS/CC/SCALbx10_ARA0 te=63-te-63 write args=0, 11, C16(97);@16_SS/CC/SCALbx14_ARC0 te=63-te-63 write args=0, 13, C16(101)                                                                                                                                                                                                                                         |
| 64  | 900 | W64 DATA  | @_UINT/CC/SCALbx34_ARA0 te=64-te-64 write args=0, 191, Cu(-2056179517);@_SINT/CC/SCALbx16_ARA0 te=64-te-64 write args=0, 335, C(1);@16_SS/CC/SCALbx10_ARA0 te=64-te-64 write args=0, 10, C16(121);@16_SS/CC/SCALbx14_ARC0 te=64-te-64 write args=0, 12, C16(113)                                                                                                                                                                                                                                       |
| 65  | 900 | W65 DATA  | @_UINT/CC/SCALbx34_ARA0 te=65-te-65 write args=0, 190, Cu(-2119160460);@_SINT/CC/SCALbx16_ARA0 te=65-te-65 write args=0, 334, C(-1);@16_SS/CC/SCALbx10_ARA0 te=65-te-65 write args=0, 9, C16(101);@16_SS/CC/SCALbx14_ARC0 te=65-te-65 write args=0, 11, C16(107)                                                                                                                                                                                                                                       |
| 66  | 900 | W66 DATA  | @_UINT/CC/SCALbx34_ARA0 te=66-te-66 write args=0, 189, Cu(-1930228819);@_SINT/CC/SCALbx16_ARA0 te=66-te-66 write args=0, 333, C(-1);@16_SS/CC/SCALbx10_ARA0 te=66-te-66 write args=0, 8, C16(112);@16_SS/CC/SCALbx14_ARC0 te=66-te-66 write args=0, 10, C16(97)                                                                                                                                                                                                                                        |
| 67  | 900 | W67 DATA  | @_UINT/CC/SCALbx34_ARA0 te=67-te-67 write args=0, 188, Cu(-2009983462);@_SINT/CC/SCALbx16_ARA0 te=67-te-67 write args=0, 332, C(0);@16_SS/CC/SCALbx10_ARA0 te=67-te-67 write args=0, 7, C16(114);@16_SS/CC/SCALbx14_ARC0 te=67-te-67 write args=0, 9, C16(101)                                                                                                                                                                                                                                         |
| 68  | 900 | W68 DATA  | @_UINT/CC/SCALbx34_ARA0 te=68-te-68 write args=0, 187, Cu(-1770699233);@_SINT/CC/SCALbx16_ARA0 te=68-te-68 write args=0, 331, C(0);@16_SS/CC/SCALbx10_ARA0 te=68-te-68 write args=0, 6, C16(102);@16_SS/CC/SCALbx14_ARC0 te=68-te-68 write args=0, 8, C16(116)                                                                                                                                                                                                                                         |
| 69  | 900 | W69 DATA  | @_UINT/CC/SCALbx34_ARA0 te=69-te-69 write args=0, 186, Cu(-1833673816);@_SINT/CC/SCALbx16_ARA0 te=69-te-69 write args=0, 330, C(-1);@16_SS/CC/SCALbx10_ARA0 te=69-te-69 write args=0, 5, C16(112);@16_SS/CC/SCALbx14_ARC0 te=69-te-69 write args=0, 7, C16(107)                                                                                                                                                                                                                                        |
| 70  | 900 | W70 DATA  | @_UINT/CC/SCALbx34_ARA0 te=70-te-70 write args=0, 185, Cu(-1611170447);@_SINT/CC/SCALbx16_ARA0 te=70-te-70 write args=0, 329, C(-2);@16_SS/CC/SCALbx10_ARA0 te=70-te-70 write args=0, 4, C16(105);@16_SS/CC/SCALbx14_ARC0 te=70-te-70 write args=0, 6, C16(116)                                                                                                                                                                                                                                        |
| 71  | 900 | W71 DATA  | @_UINT/CC/SCALbx34_ARA0 te=71-te-71 write args=0, 184, Cu(-1690935098);@_SINT/CC/SCALbx16_ARA0 te=71-te-71 write args=0, 328, C(0);@16_SS/CC/SCALbx10_ARA0 te=71-te-71 write args=0, 3, C16(97);@16_SS/CC/SCALbx14_ARC0 te=71-te-71 write args=0, 5, C16(105)                                                                                                                                                                                                                                          |
| 72  | 900 | W72 DATA  | @_UINT/CC/SCALbx34_ARA0 te=72-te-72 write args=0, 183, Cu(-1552294533);@_SINT/CC/SCALbx16_ARA0 te=72-te-72 write args=0, 327, C(0);@16_SS/CC/SCALbx10_ARA0 te=72-te-72 write args=0, 2, C16(101);@16_SS/CC/SCALbx14_ARC0 te=72-te-72 write args=0, 4, C16(108)                                                                                                                                                                                                                                         |
| 73  | 900 | W73 DATA  | @_UINT/CC/SCALbx34_ARA0 te=73-te-73 write args=0, 182, Cu(-1481064244);@_SINT/CC/SCALbx16_ARA0 te=73-te-73 write args=0, 326, C(-1);@16_SS/CC/SCALbx10_ARA0 te=73-te-73 write args=0, 1, C16(112);@16_SS/CC/SCALbx14_ARC0 te=73-te-73 write args=0, 3, C16(107)                                                                                                                                                                                                                                        |
| 74  | 900 | W74 DATA  | @_UINT/CC/SCALbx34_ARA0 te=74-te-74 write args=0, 181, Cu(-1426332139);@_SINT/CC/SCALbx16_ARA0 te=74-te-74 write args=0, 325, C(0);@16_SS/CC/SCALbx10_ARA0 te=74-te-74 write args=0, 0, C16(112);@16_SS/CC/SCALbx14_ARC0 te=74-te-74 write args=0, 2, C16(104)                                                                                                                                                                                                                                         |
| 75  | 900 | W75 DATA  | @_UINT/CC/SCALbx34_ARA0 te=75-te-75 write args=0, 180, Cu(-1371866206);@_SINT/CC/SCALbx16_ARA0 te=75-te-75 write args=0, 324, C(-3);@16_SS/CC/SCALbx14_ARC0 te=75-te-75 write args=0, 1, C16(107)                                                                                                                                                                                                                                                                                                      |
| 76  | 900 | W76 DATA  | @_UINT/CC/SCALbx34_ARA0 te=76-te-76 write args=0, 179, Cu(-1333941337);@_SINT/CC/SCALbx16_ARA0 te=76-te-76 write args=0, 323, C(0);@16_SS/CC/SCALbx14_ARC0 te=76-te-76 write args=0, 0, C16(100)                                                                                                                                                                                                                                                                                                       |
| 77  | 900 | W77 DATA  | @_UINT/CC/SCALbx34_ARA0 te=77-te-77 write args=0, 178, Cu(-1262701040);@_SINT/CC/SCALbx16_ARA0 te=77-te-77 write args=0, 322, C(0)                                                                                                                                                                                                                                                                                                                                                                     |
| 78  | 900 | W78 DATA  | @_UINT/CC/SCALbx34_ARA0 te=78-te-78 write args=0, 177, Cu(-1174433591);@_SINT/CC/SCALbx16_ARA0 te=78-te-78 write args=0, 321, C(-2)                                                                                                                                                                                                                                                                                                                                                                    |
| 79  | 900 | W79 DATA  | @_UINT/CC/SCALbx34_ARA0 te=79-te-79 write args=0, 176, Cu(-1119974018);@_SINT/CC/SCALbx16_ARA0 te=79-te-79 write args=0, 320, C(1)                                                                                                                                                                                                                                                                                                                                                                     |
| 80  | 900 | W80 DATA  | @_UINT/CC/SCALbx34_ARA0 te=80-te-80 write args=0, 175, Cu(-916395085);@_SINT/CC/SCALbx16_ARA0 te=80-te-80 write args=0, 319, C(-3)                                                                                                                                                                                                                                                                                                                                                                     |
| 81  | 900 | W81 DATA  | @_UINT/CC/SCALbx34_ARA0 te=81-te-81 write args=0, 174, Cu(-845023740);@_SINT/CC/SCALbx16_ARA0 te=81-te-81 write args=0, 318, C(-2)                                                                                                                                                                                                                                                                                                                                                                     |
| 82  | 900 | W82 DATA  | @_UINT/CC/SCALbx34_ARA0 te=82-te-82 write args=0, 173, Cu(-1058877219);@_SINT/CC/SCALbx16_ARA0 te=82-te-82 write args=0, 317, C(-1)                                                                                                                                                                                                                                                                                                                                                                    |
| 83  | 900 | W83 DATA  | @_UINT/CC/SCALbx34_ARA0 te=83-te-83 write args=0, 172, Cu(-1004286614);@_SINT/CC/SCALbx16_ARA0 te=83-te-83 write args=0, 316, C(1)                                                                                                                                                                                                                                                                                                                                                                     |
| 84  | 900 | W84 DATA  | @_UINT/CC/SCALbx34_ARA0 te=84-te-84 write args=0, 171, Cu(-630940305);@_SINT/CC/SCALbx16_ARA0 te=84-te-84 write args=0, 315, C(2)                                                                                                                                                                                                                                                                                                                                                                      |
| 85  | 900 | W85 DATA  | @_UINT/CC/SCALbx34_ARA0 te=85-te-85 write args=0, 170, Cu(-559578920);@_SINT/CC/SCALbx16_ARA0 te=85-te-85 write args=0, 314, C(0)                                                                                                                                                                                                                                                                                                                                                                      |
| 86  | 900 | W86 DATA  | @_UINT/CC/SCALbx34_ARA0 te=86-te-86 write args=0, 169, Cu(-739858943);@_SINT/CC/SCALbx16_ARA0 te=86-te-86 write args=0, 313, C(-1)                                                                                                                                                                                                                                                                                                                                                                     |
| 87  | 900 | W87 DATA  | @_UINT/CC/SCALbx34_ARA0 te=87-te-87 write args=0, 168, Cu(-685261898);@_SINT/CC/SCALbx16_ARA0 te=87-te-87 write args=0, 312, C(1)                                                                                                                                                                                                                                                                                                                                                                      |
| 88  | 900 | W88 DATA  | @_UINT/CC/SCALbx34_ARA0 te=88-te-88 write args=0, 167, Cu(-278395381);@_SINT/CC/SCALbx16_ARA0 te=88-te-88 write args=0, 311, C(1)                                                                                                                                                                                                                                                                                                                                                                      |
| 89  | 900 | W89 DATA  | @_UINT/CC/SCALbx34_ARA0 te=89-te-89 write args=0, 166, Cu(-341238852);@_SINT/CC/SCALbx16_ARA0 te=89-te-89 write args=0, 310, C(-2)                                                                                                                                                                                                                                                                                                                                                                     |
| 90  | 900 | W90 DATA  | @_UINT/CC/SCALbx34_ARA0 te=90-te-90 write args=0, 165, Cu(-420856475);@_SINT/CC/SCALbx16_ARA0 te=90-te-90 write args=0, 309, C(-3)                                                                                                                                                                                                                                                                                                                                                                     |
| 91  | 900 | W91 DATA  | @_UINT/CC/SCALbx34_ARA0 te=91-te-91 write args=0, 164, Cu(-500490030);@_SINT/CC/SCALbx16_ARA0 te=91-te-91 write args=0, 308, C(0)                                                                                                                                                                                                                                                                                                                                                                      |
| 92  | 900 | W92 DATA  | @_UINT/CC/SCALbx34_ARA0 te=92-te-92 write args=0, 163, Cu(-60002089);@_SINT/CC/SCALbx16_ARA0 te=92-te-92 write args=0, 307, C(-1)                                                                                                                                                                                                                                                                                                                                                                      |
| 93  | 900 | W93 DATA  | @_UINT/CC/SCALbx34_ARA0 te=93-te-93 write args=0, 162, Cu(-122852000);@_SINT/CC/SCALbx16_ARA0 te=93-te-93 write args=0, 306, C(-1)                                                                                                                                                                                                                                                                                                                                                                     |
| 94  | 900 | W94 DATA  | @_UINT/CC/SCALbx34_ARA0 te=94-te-94 write args=0, 161, Cu(-168932423);@_SINT/CC/SCALbx16_ARA0 te=94-te-94 write args=0, 305, C(1)                                                                                                                                                                                                                                                                                                                                                                      |
| 95  | 900 | W95 DATA  | @_UINT/CC/SCALbx34_ARA0 te=95-te-95 write args=0, 160, Cu(-248556018);@_SINT/CC/SCALbx16_ARA0 te=95-te-95 write args=0, 304, C(-3)                                                                                                                                                                                                                                                                                                                                                                     |
| 96  | 900 | W96 DATA  | @_UINT/CC/SCALbx34_ARA0 te=96-te-96 write args=0, 159, Cu(491947555);@_SINT/CC/SCALbx16_ARA0 te=96-te-96 write args=0, 303, C(0)                                                                                                                                                                                                                                                                                                                                                                       |
| 97  | 900 | W97 DATA  | @_UINT/CC/SCALbx34_ARA0 te=97-te-97 write args=0, 158, Cu(429104020);@_SINT/CC/SCALbx16_ARA0 te=97-te-97 write args=0, 302, C(0)                                                                                                                                                                                                                                                                                                                                                                       |
| 98  | 900 | W98 DATA  | @_UINT/CC/SCALbx34_ARA0 te=98-te-98 write args=0, 157, Cu(349224269);@_SINT/CC/SCALbx16_ARA0 te=98-te-98 write args=0, 301, C(0)                                                                                                                                                                                                                                                                                                                                                                       |
| 99  | 900 | W99 DATA  | @_UINT/CC/SCALbx34_ARA0 te=99-te-99 write args=0, 156, Cu(269590778);@_SINT/CC/SCALbx16_ARA0 te=99-te-99 write args=0, 300, C(1)                                                                                                                                                                                                                                                                                                                                                                       |
| 100 | 900 | W100 DATA | @_UINT/CC/SCALbx34_ARA0 te=100-te-100 write args=0, 155, Cu(240578815);@_SINT/CC/SCALbx16_ARA0 te=100-te-100 write args=0, 299, C(-4)                                                                                                                                                                                                                                                                                                                                                                  |
| 101 | 900 | W101 DATA | @_UINT/CC/SCALbx34_ARA0 te=101-te-101 write args=0, 154, Cu(177728840);@_SINT/CC/SCALbx16_ARA0 te=101-te-101 write args=0, 298, C(2)                                                                                                                                                                                                                                                                                                                                                                   |
| 102 | 900 | W102 DATA | @_UINT/CC/SCALbx34_ARA0 te=102-te-102 write args=0, 153, Cu(131386257);@_SINT/CC/SCALbx16_ARA0 te=102-te-102 write args=0, 297, C(-2)                                                                                                                                                                                                                                                                                                                                                                  |
| 103 | 900 | W103 DATA | @_UINT/CC/SCALbx34_ARA0 te=103-te-103 write args=0, 152, Cu(51762726);@_SINT/CC/SCALbx16_ARA0 te=103-te-103 write args=0, 296, C(-1)                                                                                                                                                                                                                                                                                                                                                                   |
| 104 | 900 | W104 DATA | @_UINT/CC/SCALbx34_ARA0 te=104-te-104 write args=0, 151, Cu(995781531);@_SINT/CC/SCALbx16_ARA0 te=104-te-104 write args=0, 295, C(0)                                                                                                                                                                                                                                                                                                                                                                   |
| 105 | 900 | W105 DATA | @_UINT/CC/SCALbx34_ARA0 te=105-te-105 write args=0, 150, Cu(1067152940);@_SINT/CC/SCALbx16_ARA0 te=105-te-105 write args=0, 294, C(6)                                                                                                                                                                                                                                                                                                                                                                  |
| 106 | 900 | W106 DATA | @_UINT/CC/SCALbx34_ARA0 te=106-te-106 write args=0, 149, Cu(853037301);@_SINT/CC/SCALbx16_ARA0 te=106-te-106 write args=0, 293, C(1)                                                                                                                                                                                                                                                                                                                                                                   |
| 107 | 900 | W107 DATA | @_UINT/CC/SCALbx34_ARA0 te=107-te-107 write args=0, 148, Cu(907627842);@_SINT/CC/SCALbx16_ARA0 te=107-te-107 write args=0, 292, C(0)                                                                                                                                                                                                                                                                                                                                                                   |
| 108 | 900 | W108 DATA | @_UINT/CC/SCALbx34_ARA0 te=108-te-108 write args=0, 147, Cu(677256519);@_SINT/CC/SCALbx16_ARA0 te=108-te-108 write args=0, 291, C(0)                                                                                                                                                                                                                                                                                                                                                                   |
| 109 | 900 | W109 DATA | @_UINT/CC/SCALbx34_ARA0 te=109-te-109 write args=0, 146, Cu(748617968);@_SINT/CC/SCALbx16_ARA0 te=109-te-109 write args=0, 290, C(0)                                                                                                                                                                                                                                                                                                                                                                   |
| 110 | 900 | W110 DATA | @_UINT/CC/SCALbx34_ARA0 te=110-te-110 write args=0, 145, Cu(568075817);@_SINT/CC/SCALbx16_ARA0 te=110-te-110 write args=0, 289, C(-3)                                                                                                                                                                                                                                                                                                                                                                  |
| 111 | 900 | W111 DATA | @_UINT/CC/SCALbx34_ARA0 te=111-te-111 write args=0, 144, Cu(622672798);@_SINT/CC/SCALbx16_ARA0 te=111-te-111 write args=0, 288, C(3)                                                                                                                                                                                                                                                                                                                                                                   |
| 112 | 900 | W112 DATA | @_UINT/CC/SCALbx34_ARA0 te=112-te-112 write args=0, 143, Cu(1363369299);@_SINT/CC/SCALbx16_ARA0 te=112-te-112 write args=0, 287, C(-2)                                                                                                                                                                                                                                                                                                                                                                 |
| 113 | 900 | W113 DATA | @_UINT/CC/SCALbx34_ARA0 te=113-te-113 write args=0, 142, Cu(1434599652);@_SINT/CC/SCALbx16_ARA0 te=113-te-113 write args=0, 286, C(2)                                                                                                                                                                                                                                                                                                                                                                  |
| 114 | 900 | W114 DATA | @_UINT/CC/SCALbx34_ARA0 te=114-te-114 write args=0, 141, Cu(1489069629);@_SINT/CC/SCALbx16_ARA0 te=114-te-114 write args=0, 285, C(-3)                                                                                                                                                                                                                                                                                                                                                                 |
| 115 | 900 | W115 DATA | @_UINT/CC/SCALbx34_ARA0 te=115-te-115 write args=0, 140, Cu(1543535498);@_SINT/CC/SCALbx16_ARA0 te=115-te-115 write args=0, 284, C(-4)                                                                                                                                                                                                                                                                                                                                                                 |
| 116 | 900 | W116 DATA | @_UINT/CC/SCALbx34_ARA0 te=116-te-116 write args=0, 139, Cu(1111960463);@_SINT/CC/SCALbx16_ARA0 te=116-te-116 write args=0, 283, C(-1)                                                                                                                                                                                                                                                                                                                                                                 |
| 117 | 900 | W117 DATA | @_UINT/CC/SCALbx34_ARA0 te=117-te-117 write args=0, 138, Cu(1183200824);@_SINT/CC/SCALbx16_ARA0 te=117-te-117 write args=0, 282, C(-1)                                                                                                                                                                                                                                                                                                                                                                 |
| 118 | 900 | W118 DATA | @_UINT/CC/SCALbx34_ARA0 te=118-te-118 write args=0, 137, Cu(1271206113);@_SINT/CC/SCALbx16_ARA0 te=118-te-118 write args=0, 281, C(-4)                                                                                                                                                                                                                                                                                                                                                                 |
| 119 | 900 | W119 DATA | @_UINT/CC/SCALbx34_ARA0 te=119-te-119 write args=0, 136, Cu(1325665622);@_SINT/CC/SCALbx16_ARA0 te=119-te-119 write args=0, 280, C(-2)                                                                                                                                                                                                                                                                                                                                                                 |
| 120 | 900 | W120 DATA | @_UINT/CC/SCALbx34_ARA0 te=120-te-120 write args=0, 135, Cu(2001449195);@_SINT/CC/SCALbx16_ARA0 te=120-te-120 write args=0, 279, C(-4)                                                                                                                                                                                                                                                                                                                                                                 |
| 121 | 900 | W121 DATA | @_UINT/CC/SCALbx34_ARA0 te=121-te-121 write args=0, 134, Cu(1938468188);@_SINT/CC/SCALbx16_ARA0 te=121-te-121 write args=0, 278, C(-5)                                                                                                                                                                                                                                                                                                                                                                 |
| 122 | 900 | W122 DATA | @_UINT/CC/SCALbx34_ARA0 te=122-te-122 write args=0, 133, Cu(2127137669);@_SINT/CC/SCALbx16_ARA0 te=122-te-122 write args=0, 277, C(-2)                                                                                                                                                                                                                                                                                                                                                                 |
| 123 | 900 | W123 DATA | @_UINT/CC/SCALbx34_ARA0 te=123-te-123 write args=0, 132, Cu(2047383090);@_SINT/CC/SCALbx16_ARA0 te=123-te-123 write args=0, 276, C(-1)                                                                                                                                                                                                                                                                                                                                                                 |
| 124 | 900 | W124 DATA | @_UINT/CC/SCALbx34_ARA0 te=124-te-124 write args=0, 131, Cu(1682949687);@_SINT/CC/SCALbx16_ARA0 te=124-te-124 write args=0, 275, C(-1)                                                                                                                                                                                                                                                                                                                                                                 |
| 125 | 900 | W125 DATA | @_UINT/CC/SCALbx34_ARA0 te=125-te-125 write args=0, 130, Cu(1619975040);@_SINT/CC/SCALbx16_ARA0 te=125-te-125 write args=0, 274, C(1)                                                                                                                                                                                                                                                                                                                                                                  |
| 126 | 900 | W126 DATA | @_UINT/CC/SCALbx34_ARA0 te=126-te-126 write args=0, 129, Cu(1842216281);@_SINT/CC/SCALbx16_ARA0 te=126-te-126 write args=0, 273, C(4)                                                                                                                                                                                                                                                                                                                                                                  |
| 127 | 900 | W127 DATA | @_UINT/CC/SCALbx34_ARA0 te=127-te-127 write args=0, 128, Cu(1762451694);@_SINT/CC/SCALbx16_ARA0 te=127-te-127 write args=0, 272, C(0)                                                                                                                                                                                                                                                                                                                                                                  |
| 128 | 900 | W128 DATA | @_UINT/CC/SCALbx34_ARA0 te=128-te-128 write args=0, 127, Cu(-654598054);@_SINT/CC/SCALbx16_ARA0 te=128-te-128 write args=0, 271, C(1)                                                                                                                                                                                                                                                                                                                                                                  |
| 129 | 900 | W129 DATA | @_UINT/CC/SCALbx34_ARA0 te=129-te-129 write args=0, 126, Cu(-600130067);@_SINT/CC/SCALbx16_ARA0 te=129-te-129 write args=0, 270, C(-1)                                                                                                                                                                                                                                                                                                                                                                 |
| 130 | 900 | W130 DATA | @_UINT/CC/SCALbx34_ARA0 te=130-te-130 write args=0, 125, Cu(-780559564);@_SINT/CC/SCALbx16_ARA0 te=130-te-130 write args=0, 269, C(-2)                                                                                                                                                                                                                                                                                                                                                                 |
| 131 | 900 | W131 DATA | @_UINT/CC/SCALbx34_ARA0 te=131-te-131 write args=0, 124, Cu(-709327229);@_SINT/CC/SCALbx16_ARA0 te=131-te-131 write args=0, 268, C(1)                                                                                                                                                                                                                                                                                                                                                                  |
| 132 | 900 | W132 DATA | @_UINT/CC/SCALbx34_ARA0 te=132-te-132 write args=0, 123, Cu(-872425850);@_SINT/CC/SCALbx16_ARA0 te=132-te-132 write args=0, 267, C(-2)                                                                                                                                                                                                                                                                                                                                                                 |
| 133 | 900 | W133 DATA | @_UINT/CC/SCALbx34_ARA0 te=133-te-133 write args=0, 122, Cu(-817968335);@_SINT/CC/SCALbx16_ARA0 te=133-te-133 write args=0, 266, C(3)                                                                                                                                                                                                                                                                                                                                                                  |
| 134 | 900 | W134 DATA | @_UINT/CC/SCALbx34_ARA0 te=134-te-134 write args=0, 121, Cu(-1031934488);@_SINT/CC/SCALbx16_ARA0 te=134-te-134 write args=0, 265, C(-1)                                                                                                                                                                                                                                                                                                                                                                |
| 135 | 900 | W135 DATA | @_UINT/CC/SCALbx34_ARA0 te=135-te-135 write args=0, 120, Cu(-960696225);@_SINT/CC/SCALbx16_ARA0 te=135-te-135 write args=0, 264, C(-5)                                                                                                                                                                                                                                                                                                                                                                 |
| 136 | 900 | W136 DATA | @_UINT/CC/SCALbx34_ARA0 te=136-te-136 write args=0, 119, Cu(-17609246);@_SINT/CC/SCALbx16_ARA0 te=136-te-136 write args=0, 263, C(2)                                                                                                                                                                                                                                                                                                                                                                   |
| 137 | 900 | W137 DATA | @_UINT/CC/SCALbx34_ARA0 te=137-te-137 write args=0, 118, Cu(-97365931);@_SINT/CC/SCALbx16_ARA0 te=137-te-137 write args=0, 262, C(2)                                                                                                                                                                                                                                                                                                                                                                   |
| 138 | 900 | W138 DATA | @_UINT/CC/SCALbx34_ARA0 te=138-te-138 write args=0, 117, Cu(-143559028);@_SINT/CC/SCALbx16_ARA0 te=138-te-138 write args=0, 261, C(-5)                                                                                                                                                                                                                                                                                                                                                                 |
| 139 | 900 | W139 DATA | @_UINT/CC/SCALbx34_ARA0 te=139-te-139 write args=0, 116, Cu(-206542021);@_SINT/CC/SCALbx16_ARA0 te=139-te-139 write args=0, 260, C(0)                                                                                                                                                                                                                                                                                                                                                                  |
| 140 | 900 | W140 DATA | @_UINT/CC/SCALbx34_ARA0 te=140-te-140 write args=0, 115, Cu(-302564546);@_SINT/CC/SCALbx16_ARA0 te=140-te-140 write args=0, 259, C(-5)                                                                                                                                                                                                                                                                                                                                                                 |
| 141 | 900 | W141 DATA | @_UINT/CC/SCALbx34_ARA0 te=141-te-141 write args=0, 114, Cu(-382327159);@_SINT/CC/SCALbx16_ARA0 te=141-te-141 write args=0, 258, C(-6)                                                                                                                                                                                                                                                                                                                                                                 |
| 142 | 900 | W142 DATA | @_UINT/CC/SCALbx34_ARA0 te=142-te-142 write args=0, 113, Cu(-462094256);@_SINT/CC/SCALbx16_ARA0 te=142-te-142 write args=0, 257, C(-1)                                                                                                                                                                                                                                                                                                                                                                 |
| 143 | 900 | W143 DATA | @_UINT/CC/SCALbx34_ARA0 te=143-te-143 write args=0, 112, Cu(-525066777);@_SINT/CC/SCALbx16_ARA0 te=143-te-143 write args=0, 256, C(0)                                                                                                                                                                                                                                                                                                                                                                  |
| 144 | 900 | W144 DATA | @_UINT/CC/SCALbx34_ARA0 te=144-te-144 write args=0, 111, Cu(-1796572374);@_SINT/CC/SCALbx16_ARA0 te=144-te-144 write args=0, 255, C(1)                                                                                                                                                                                                                                                                                                                                                                 |
| 145 | 900 | W145 DATA | @_UINT/CC/SCALbx34_ARA0 te=145-te-145 write args=0, 110, Cu(-1876203875);@_SINT/CC/SCALbx16_ARA0 te=145-te-145 write args=0, 254, C(0)                                                                                                                                                                                                                                                                                                                                                                 |
| 146 | 900 | W146 DATA | @_UINT/CC/SCALbx34_ARA0 te=146-te-146 write args=0, 109, Cu(-1654112188);@_SINT/CC/SCALbx16_ARA0 te=146-te-146 write args=0, 253, C(0)                                                                                                                                                                                                                                                                                                                                                                 |
| 147 | 900 | W147 DATA | @_UINT/CC/SCALbx34_ARA0 te=147-te-147 write args=0, 108, Cu(-1716953613);@_SINT/CC/SCALbx16_ARA0 te=147-te-147 write args=0, 252, C(6)                                                                                                                                                                                                                                                                                                                                                                 |
| 148 | 900 | W148 DATA | @_UINT/CC/SCALbx34_ARA0 te=148-te-148 write args=0, 107, Cu(-2014441994);@_SINT/CC/SCALbx16_ARA0 te=148-te-148 write args=0, 251, C(-1)                                                                                                                                                                                                                                                                                                                                                                |
| 149 | 900 | W149 DATA | @_UINT/CC/SCALbx34_ARA0 te=149-te-149 write args=0, 106, Cu(-2094067647);@_SINT/CC/SCALbx16_ARA0 te=149-te-149 write args=0, 250, C(-2)                                                                                                                                                                                                                                                                                                                                                                |
| 150 | 900 | W150 DATA | @_UINT/CC/SCALbx34_ARA0 te=150-te-150 write args=0, 105, Cu(-1905510760);@_SINT/CC/SCALbx16_ARA0 te=150-te-150 write args=0, 249, C(-3)                                                                                                                                                                                                                                                                                                                                                                |
| 151 | 900 | W151 DATA | @_UINT/CC/SCALbx34_ARA0 te=151-te-151 write args=0, 104, Cu(-1968362705);@_SINT/CC/SCALbx16_ARA0 te=151-te-151 write args=0, 248, C(-1)                                                                                                                                                                                                                                                                                                                                                                |
| 152 | 900 | W152 DATA | @_UINT/CC/SCALbx34_ARA0 te=152-te-152 write args=0, 103, Cu(-1293773166);@_SINT/CC/SCALbx16_ARA0 te=152-te-152 write args=0, 247, C(-2)                                                                                                                                                                                                                                                                                                                                                                |
| 153 | 900 | W153 DATA | @_UINT/CC/SCALbx34_ARA0 te=153-te-153 write args=0, 102, Cu(-1239184603);@_SINT/CC/SCALbx16_ARA0 te=153-te-153 write args=0, 246, C(0)                                                                                                                                                                                                                                                                                                                                                                 |
| 154 | 900 | W154 DATA | @_UINT/CC/SCALbx34_ARA0 te=154-te-154 write args=0, 101, Cu(-1151291908);@_SINT/CC/SCALbx16_ARA0 te=154-te-154 write args=0, 245, C(-1)                                                                                                                                                                                                                                                                                                                                                                |
| 155 | 900 | W155 DATA | @_UINT/CC/SCALbx34_ARA0 te=155-te-155 write args=0, 100, Cu(-1079922613);@_SINT/CC/SCALbx16_ARA0 te=155-te-155 write args=0, 244, C(-5)                                                                                                                                                                                                                                                                                                                                                                |
| 156 | 900 | W156 DATA | @_UINT/CC/SCALbx34_ARA0 te=156-te-156 write args=0, 99, Cu(-1578704818);@_SINT/CC/SCALbx16_ARA0 te=156-te-156 write args=0, 243, C(-1)                                                                                                                                                                                                                                                                                                                                                                 |
| 157 | 900 | W157 DATA | @_UINT/CC/SCALbx34_ARA0 te=157-te-157 write args=0, 98, Cu(-1524105735);@_SINT/CC/SCALbx16_ARA0 te=157-te-157 write args=0, 242, C(-1)                                                                                                                                                                                                                                                                                                                                                                 |
| 158 | 900 | W158 DATA | @_UINT/CC/SCALbx34_ARA0 te=158-te-158 write args=0, 97, Cu(-1469785312);@_SINT/CC/SCALbx16_ARA0 te=158-te-158 write args=0, 241, C(-3)                                                                                                                                                                                                                                                                                                                                                                 |
| 159 | 900 | W159 DATA | @_UINT/CC/SCALbx34_ARA0 te=159-te-159 write args=0, 96, Cu(-1398421865);@_SINT/CC/SCALbx16_ARA0 te=159-te-159 write args=0, 240, C(1)                                                                                                                                                                                                                                                                                                                                                                  |
| 160 | 900 | W160 DATA | @_UINT/CC/SCALbx34_ARA0 te=160-te-160 write args=0, 95, Cu(1087903418);@_SINT/CC/SCALbx16_ARA0 te=160-te-160 write args=0, 239, C(-2)                                                                                                                                                                                                                                                                                                                                                                  |
| 161 | 900 | W161 DATA | @_UINT/CC/SCALbx34_ARA0 te=161-te-161 write args=0, 94, Cu(1142491917);@_SINT/CC/SCALbx16_ARA0 te=161-te-161 write args=0, 238, C(-4)                                                                                                                                                                                                                                                                                                                                                                  |
| 162 | 900 | W162 DATA | @_UINT/CC/SCALbx34_ARA0 te=162-te-162 write args=0, 93, Cu(1230646740);@_SINT/CC/SCALbx16_ARA0 te=162-te-162 write args=0, 237, C(-2)                                                                                                                                                                                                                                                                                                                                                                  |
| 163 | 900 | W163 DATA | @_UINT/CC/SCALbx34_ARA0 te=163-te-163 write args=0, 92, Cu(1302016099);@_SINT/CC/SCALbx16_ARA0 te=163-te-163 write args=0, 236, C(0)                                                                                                                                                                                                                                                                                                                                                                   |
| 164 | 900 | W164 DATA | @_UINT/CC/SCALbx34_ARA0 te=164-te-164 write args=0, 91, Cu(1406951526);@_SINT/CC/SCALbx16_ARA0 te=164-te-164 write args=0, 235, C(1)                                                                                                                                                                                                                                                                                                                                                                   |
| 165 | 900 | W165 DATA | @_UINT/CC/SCALbx34_ARA0 te=165-te-165 write args=0, 90, Cu(1461550545);@_SINT/CC/SCALbx16_ARA0 te=165-te-165 write args=0, 234, C(0)                                                                                                                                                                                                                                                                                                                                                                   |
| 166 | 900 | W166 DATA | @_UINT/CC/SCALbx34_ARA0 te=166-te-166 write args=0, 89, Cu(1516133128);@_SINT/CC/SCALbx16_ARA0 te=166-te-166 write args=0, 233, C(1)                                                                                                                                                                                                                                                                                                                                                                   |
| 167 | 900 | W167 DATA | @_UINT/CC/SCALbx34_ARA0 te=167-te-167 write args=0, 88, Cu(1587496639);@_SINT/CC/SCALbx16_ARA0 te=167-te-167 write args=0, 232, C(-1)                                                                                                                                                                                                                                                                                                                                                                  |
| 168 | 900 | W168 DATA | @_UINT/CC/SCALbx34_ARA0 te=168-te-168 write args=0, 87, Cu(1724971778);@_SINT/CC/SCALbx16_ARA0 te=168-te-168 write args=0, 231, C(2)                                                                                                                                                                                                                                                                                                                                                                   |
| 169 | 900 | W169 DATA | @_UINT/CC/SCALbx34_ARA0 te=169-te-169 write args=0, 86, Cu(1645340341);@_SINT/CC/SCALbx16_ARA0 te=169-te-169 write args=0, 230, C(-2)                                                                                                                                                                                                                                                                                                                                                                  |
| 170 | 900 | W170 DATA | @_UINT/CC/SCALbx34_ARA0 te=170-te-170 write args=0, 85, Cu(1867694188);@_SINT/CC/SCALbx16_ARA0 te=170-te-170 write args=0, 229, C(-3)                                                                                                                                                                                                                                                                                                                                                                  |
| 171 | 900 | W171 DATA | @_UINT/CC/SCALbx34_ARA0 te=171-te-171 write args=0, 84, Cu(1804852699);@_SINT/CC/SCALbx16_ARA0 te=171-te-171 write args=0, 228, C(1)                                                                                                                                                                                                                                                                                                                                                                   |
| 172 | 900 | W172 DATA | @_UINT/CC/SCALbx34_ARA0 te=172-te-172 write args=0, 83, Cu(1976864222);@_SINT/CC/SCALbx16_ARA0 te=172-te-172 write args=0, 227, C(-2)                                                                                                                                                                                                                                                                                                                                                                  |
| 173 | 900 | W173 DATA | @_UINT/CC/SCALbx34_ARA0 te=173-te-173 write args=0, 82, Cu(1897238633);@_SINT/CC/SCALbx16_ARA0 te=173-te-173 write args=0, 226, C(2)                                                                                                                                                                                                                                                                                                                                                                   |
| 174 | 900 | W174 DATA | @_UINT/CC/SCALbx34_ARA0 te=174-te-174 write args=0, 81, Cu(2086057648);@_SINT/CC/SCALbx16_ARA0 te=174-te-174 write args=0, 225, C(0)                                                                                                                                                                                                                                                                                                                                                                   |
| 175 | 900 | W175 DATA | @_UINT/CC/SCALbx34_ARA0 te=175-te-175 write args=0, 80, Cu(2023205639);@_SINT/CC/SCALbx16_ARA0 te=175-te-175 write args=0, 224, C(-4)                                                                                                                                                                                                                                                                                                                                                                  |
| 176 | 900 | W176 DATA | @_UINT/CC/SCALbx34_ARA0 te=176-te-176 write args=0, 79, Cu(214552010);@_SINT/CC/SCALbx16_ARA0 te=176-te-176 write args=0, 223, C(1)                                                                                                                                                                                                                                                                                                                                                                    |
| 177 | 900 | W177 DATA | @_UINT/CC/SCALbx34_ARA0 te=177-te-177 write args=0, 78, Cu(134795389);@_SINT/CC/SCALbx16_ARA0 te=177-te-177 write args=0, 222, C(2)                                                                                                                                                                                                                                                                                                                                                                    |
| 178 | 900 | W178 DATA | @_UINT/CC/SCALbx34_ARA0 te=178-te-178 write args=0, 77, Cu(88864420);@_SINT/CC/SCALbx16_ARA0 te=178-te-178 write args=0, 221, C(-4)                                                                                                                                                                                                                                                                                                                                                                    |
| 179 | 900 | W179 DATA | @_UINT/CC/SCALbx34_ARA0 te=179-te-179 write args=0, 76, Cu(25881363);@_SINT/CC/SCALbx16_ARA0 te=179-te-179 write args=0, 220, C(0)                                                                                                                                                                                                                                                                                                                                                                     |
| 180 | 900 | W180 DATA | @_UINT/CC/SCALbx34_ARA0 te=180-te-180 write args=0, 75, Cu(533576470);@_SINT/CC/SCALbx16_ARA0 te=180-te-180 write args=0, 219, C(-2)                                                                                                                                                                                                                                                                                                                                                                   |
| 181 | 900 | W181 DATA | @_UINT/CC/SCALbx34_ARA0 te=181-te-181 write args=0, 74, Cu(453813921);@_SINT/CC/SCALbx16_ARA0 te=181-te-181 write args=0, 218, C(-4)                                                                                                                                                                                                                                                                                                                                                                   |
| 182 | 900 | W182 DATA | @_UINT/CC/SCALbx34_ARA0 te=182-te-182 write args=0, 73, Cu(374308984);@_SINT/CC/SCALbx16_ARA0 te=182-te-182 write args=0, 217, C(2)                                                                                                                                                                                                                                                                                                                                                                    |
| 183 | 900 | W183 DATA | @_UINT/CC/SCALbx34_ARA0 te=183-te-183 write args=0, 72, Cu(311336399);@_SINT/CC/SCALbx16_ARA0 te=183-te-183 write args=0, 216, C(-1)                                                                                                                                                                                                                                                                                                                                                                   |
| 184 | 900 | W184 DATA | @_UINT/CC/SCALbx34_ARA0 te=184-te-184 write args=0, 71, Cu(717299826);@_SINT/CC/SCALbx16_ARA0 te=184-te-184 write args=0, 215, C(-2)                                                                                                                                                                                                                                                                                                                                                                   |
| 185 | 900 | W185 DATA | @_UINT/CC/SCALbx34_ARA0 te=185-te-185 write args=0, 70, Cu(771767749);@_SINT/CC/SCALbx16_ARA0 te=185-te-185 write args=0, 214, C(0)                                                                                                                                                                                                                                                                                                                                                                    |
| 186 | 900 | W186 DATA | @_UINT/CC/SCALbx34_ARA0 te=186-te-186 write args=0, 69, Cu(591600412);@_SINT/CC/SCALbx16_ARA0 te=186-te-186 write args=0, 213, C(-1)                                                                                                                                                                                                                                                                                                                                                                   |
| 187 | 900 | W187 DATA | @_UINT/CC/SCALbx34_ARA0 te=187-te-187 write args=0, 68, Cu(662832811);@_SINT/CC/SCALbx16_ARA0 te=187-te-187 write args=0, 212, C(-2)                                                                                                                                                                                                                                                                                                                                                                   |
| 188 | 900 | W188 DATA | @_UINT/CC/SCALbx34_ARA0 te=188-te-188 write args=0, 67, Cu(969234094);@_SINT/CC/SCALbx16_ARA0 te=188-te-188 write args=0, 211, C(-2)                                                                                                                                                                                                                                                                                                                                                                   |
| 189 | 900 | W189 DATA | @_UINT/CC/SCALbx34_ARA0 te=189-te-189 write args=0, 66, Cu(1023691545);@_SINT/CC/SCALbx16_ARA0 te=189-te-189 write args=0, 210, C(6)                                                                                                                                                                                                                                                                                                                                                                   |
| 190 | 900 | W190 DATA | @_UINT/CC/SCALbx34_ARA0 te=190-te-190 write args=0, 65, Cu(809987520);@_SINT/CC/SCALbx16_ARA0 te=190-te-190 write args=0, 209, C(4)                                                                                                                                                                                                                                                                                                                                                                    |
| 191 | 900 | W191 DATA | @_UINT/CC/SCALbx34_ARA0 te=191-te-191 write args=0, 64, Cu(881225847);@_SINT/CC/SCALbx16_ARA0 te=191-te-191 write args=0, 208, C(0)                                                                                                                                                                                                                                                                                                                                                                    |
| 192 | 900 | W192 DATA | @_UINT/CC/SCALbx34_ARA0 te=192-te-192 write args=0, 63, Cu(-327299027);@_SINT/CC/SCALbx16_ARA0 te=192-te-192 write args=0, 207, C(2)                                                                                                                                                                                                                                                                                                                                                                   |
| 193 | 900 | W193 DATA | @_UINT/CC/SCALbx34_ARA0 te=193-te-193 write args=0, 62, Cu(-390279782);@_SINT/CC/SCALbx16_ARA0 te=193-te-193 write args=0, 206, C(-2)                                                                                                                                                                                                                                                                                                                                                                  |
| 194 | 900 | W194 DATA | @_UINT/CC/SCALbx34_ARA0 te=194-te-194 write args=0, 61, Cu(-436212925);@_SINT/CC/SCALbx16_ARA0 te=194-te-194 write args=0, 205, C(-3)                                                                                                                                                                                                                                                                                                                                                                  |
| 195 | 900 | W195 DATA | @_UINT/CC/SCALbx34_ARA0 te=195-te-195 write args=0, 60, Cu(-515967244);@_SINT/CC/SCALbx16_ARA0 te=195-te-195 write args=0, 204, C(0)                                                                                                                                                                                                                                                                                                                                                                   |
| 196 | 900 | W196 DATA | @_UINT/CC/SCALbx34_ARA0 te=196-te-196 write args=0, 59, Cu(-8804623);@_SINT/CC/SCALbx16_ARA0 te=196-te-196 write args=0, 203, C(-2)                                                                                                                                                                                                                                                                                                                                                                    |
| 197 | 900 | W197 DATA | @_UINT/CC/SCALbx34_ARA0 te=197-te-197 write args=0, 58, Cu(-71779514);@_SINT/CC/SCALbx16_ARA0 te=197-te-197 write args=0, 202, C(-3)                                                                                                                                                                                                                                                                                                                                                                   |
| 198 | 900 | W198 DATA | @_UINT/CC/SCALbx34_ARA0 te=198-te-198 write args=0, 57, Cu(-151282273);@_SINT/CC/SCALbx16_ARA0 te=198-te-198 write args=0, 201, C(-5)                                                                                                                                                                                                                                                                                                                                                                  |
| 199 | 900 | W199 DATA | @_UINT/CC/SCALbx34_ARA0 te=199-te-199 write args=0, 56, Cu(-231047128);@_SINT/CC/SCALbx16_ARA0 te=199-te-199 write args=0, 200, C(-1)                                                                                                                                                                                                                                                                                                                                                                  |
| 200 | 900 | W200 DATA | @_UINT/CC/SCALbx34_ARA0 te=200-te-200 write args=0, 55, Cu(-898286187);@_SINT/CC/SCALbx16_ARA0 te=200-te-200 write args=0, 199, C(-1)                                                                                                                                                                                                                                                                                                                                                                  |
| 201 | 900 | W201 DATA | @_UINT/CC/SCALbx34_ARA0 te=201-te-201 write args=0, 54, Cu(-827056094);@_SINT/CC/SCALbx16_ARA0 te=201-te-201 write args=0, 198, C(-2)                                                                                                                                                                                                                                                                                                                                                                  |
| 202 | 900 | W202 DATA | @_UINT/CC/SCALbx34_ARA0 te=202-te-202 write args=0, 53, Cu(-1007220997);@_SINT/CC/SCALbx16_ARA0 te=202-te-202 write args=0, 197, C(2)                                                                                                                                                                                                                                                                                                                                                                  |
| 203 | 900 | W203 DATA | @_UINT/CC/SCALbx34_ARA0 te=203-te-203 write args=0, 52, Cu(-952755380);@_SINT/CC/SCALbx16_ARA0 te=203-te-203 write args=0, 196, C(-2)                                                                                                                                                                                                                                                                                                                                                                  |
| 204 | 900 | W204 DATA | @_UINT/CC/SCALbx34_ARA0 te=204-te-204 write args=0, 51, Cu(-646886583);@_SINT/CC/SCALbx16_ARA0 te=204-te-204 write args=0, 195, C(-3)                                                                                                                                                                                                                                                                                                                                                                  |
| 205 | 900 | W205 DATA | @_UINT/CC/SCALbx34_ARA0 te=205-te-205 write args=0, 50, Cu(-575645954);@_SINT/CC/SCALbx16_ARA0 te=205-te-205 write args=0, 194, C(-3)                                                                                                                                                                                                                                                                                                                                                                  |
| 206 | 900 | W206 DATA | @_UINT/CC/SCALbx34_ARA0 te=206-te-206 write args=0, 49, Cu(-789352409);@_SINT/CC/SCALbx16_ARA0 te=206-te-206 write args=0, 193, C(-2)                                                                                                                                                                                                                                                                                                                                                                  |
| 207 | 900 | W207 DATA | @_UINT/CC/SCALbx34_ARA0 te=207-te-207 write args=0, 48, Cu(-734892656);@_SINT/CC/SCALbx16_ARA0 te=207-te-207 write args=0, 192, C(-3)                                                                                                                                                                                                                                                                                                                                                                  |
| 208 | 900 | W208 DATA | @_UINT/CC/SCALbx34_ARA0 te=208-te-208 write args=0, 47, Cu(-1603531939);@_SINT/CC/SCALbx16_ARA0 te=208-te-208 write args=0, 191, C(-3)                                                                                                                                                                                                                                                                                                                                                                 |
| 209 | 900 | W209 DATA | @_UINT/CC/SCALbx34_ARA0 te=209-te-209 write args=0, 46, Cu(-1532160278);@_SINT/CC/SCALbx16_ARA0 te=209-te-209 write args=0, 190, C(4)                                                                                                                                                                                                                                                                                                                                                                  |
| 210 | 900 | W210 DATA | @_UINT/CC/SCALbx34_ARA0 te=210-te-210 write args=0, 45, Cu(-1444007885);@_SINT/CC/SCALbx16_ARA0 te=210-te-210 write args=0, 189, C(6)                                                                                                                                                                                                                                                                                                                                                                  |
| 211 | 900 | W211 DATA | @_UINT/CC/SCALbx34_ARA0 te=211-te-211 write args=0, 44, Cu(-1389417084);@_SINT/CC/SCALbx16_ARA0 te=211-te-211 write args=0, 188, C(-3)                                                                                                                                                                                                                                                                                                                                                                 |
| 212 | 900 | W212 DATA | @_UINT/CC/SCALbx34_ARA0 te=212-te-212 write args=0, 43, Cu(-1284997759);@_SINT/CC/SCALbx16_ARA0 te=212-te-212 write args=0, 187, C(2)                                                                                                                                                                                                                                                                                                                                                                  |
| 213 | 900 | W213 DATA | @_UINT/CC/SCALbx34_ARA0 te=213-te-213 write args=0, 42, Cu(-1213636554);@_SINT/CC/SCALbx16_ARA0 te=213-te-213 write args=0, 186, C(-2)                                                                                                                                                                                                                                                                                                                                                                 |
| 214 | 900 | W214 DATA | @_UINT/CC/SCALbx34_ARA0 te=214-te-214 write args=0, 41, Cu(-1159051537);@_SINT/CC/SCALbx16_ARA0 te=214-te-214 write args=0, 185, C(-4)                                                                                                                                                                                                                                                                                                                                                                 |
| 215 | 900 | W215 DATA | @_UINT/CC/SCALbx34_ARA0 te=215-te-215 write args=0, 40, Cu(-1104454824);@_SINT/CC/SCALbx16_ARA0 te=215-te-215 write args=0, 184, C(2)                                                                                                                                                                                                                                                                                                                                                                  |
| 216 | 900 | W216 DATA | @_UINT/CC/SCALbx34_ARA0 te=216-te-216 write args=0, 39, Cu(-2040207643);@_SINT/CC/SCALbx16_ARA0 te=216-te-216 write args=0, 183, C(-3)                                                                                                                                                                                                                                                                                                                                                                 |
| 217 | 900 | W217 DATA | @_UINT/CC/SCALbx34_ARA0 te=217-te-217 write args=0, 38, Cu(-2103051438);@_SINT/CC/SCALbx16_ARA0 te=217-te-217 write args=0, 182, C(-4)                                                                                                                                                                                                                                                                                                                                                                 |
| 218 | 900 | W218 DATA | @_UINT/CC/SCALbx34_ARA0 te=218-te-218 write args=0, 37, Cu(-1880695413);@_SINT/CC/SCALbx16_ARA0 te=218-te-218 write args=0, 181, C(-6)                                                                                                                                                                                                                                                                                                                                                                 |
| 219 | 900 | W219 DATA | @_UINT/CC/SCALbx34_ARA0 te=219-te-219 write args=0, 36, Cu(-1960329156);@_SINT/CC/SCALbx16_ARA0 te=219-te-219 write args=0, 180, C(-2)                                                                                                                                                                                                                                                                                                                                                                 |
| 220 | 900 | W220 DATA | @_UINT/CC/SCALbx34_ARA0 te=220-te-220 write args=0, 35, Cu(-1788833735);@_SINT/CC/SCALbx16_ARA0 te=220-te-220 write args=0, 179, C(-4)                                                                                                                                                                                                                                                                                                                                                                 |
| 221 | 900 | W221 DATA | @_UINT/CC/SCALbx34_ARA0 te=221-te-221 write args=0, 34, Cu(-1851683442);@_SINT/CC/SCALbx16_ARA0 te=221-te-221 write args=0, 178, C(-3)                                                                                                                                                                                                                                                                                                                                                                 |
| 222 | 900 | W222 DATA | @_UINT/CC/SCALbx34_ARA0 te=222-te-222 write args=0, 33, Cu(-1662866601);@_SINT/CC/SCALbx16_ARA0 te=222-te-222 write args=0, 177, C(-2)                                                                                                                                                                                                                                                                                                                                                                 |
| 223 | 900 | W223 DATA | @_UINT/CC/SCALbx34_ARA0 te=223-te-223 write args=0, 32, Cu(-1742489888);@_SINT/CC/SCALbx16_ARA0 te=223-te-223 write args=0, 176, C(0)                                                                                                                                                                                                                                                                                                                                                                  |
| 224 | 900 | W224 DATA | @_UINT/CC/SCALbx34_ARA0 te=224-te-224 write args=0, 31, Cu(1952343757);@_SINT/CC/SCALbx16_ARA0 te=224-te-224 write args=0, 175, C(0)                                                                                                                                                                                                                                                                                                                                                                   |
| 225 | 900 | W225 DATA | @_UINT/CC/SCALbx34_ARA0 te=225-te-225 write args=0, 30, Cu(1889500026);@_SINT/CC/SCALbx16_ARA0 te=225-te-225 write args=0, 174, C(3)                                                                                                                                                                                                                                                                                                                                                                   |
| 226 | 900 | W226 DATA | @_UINT/CC/SCALbx34_ARA0 te=226-te-226 write args=0, 29, Cu(2111593891);@_SINT/CC/SCALbx16_ARA0 te=226-te-226 write args=0, 173, C(1)                                                                                                                                                                                                                                                                                                                                                                   |
| 227 | 900 | W227 DATA | @_UINT/CC/SCALbx34_ARA0 te=227-te-227 write args=0, 28, Cu(2031960084);@_SINT/CC/SCALbx16_ARA0 te=227-te-227 write args=0, 172, C(-1)                                                                                                                                                                                                                                                                                                                                                                  |
| 228 | 900 | W228 DATA | @_UINT/CC/SCALbx34_ARA0 te=228-te-228 write args=0, 27, Cu(1733955601);@_SINT/CC/SCALbx16_ARA0 te=228-te-228 write args=0, 171, C(1)                                                                                                                                                                                                                                                                                                                                                                   |
| 229 | 900 | W229 DATA | @_UINT/CC/SCALbx34_ARA0 te=229-te-229 write args=0, 26, Cu(1671105958);@_SINT/CC/SCALbx16_ARA0 te=229-te-229 write args=0, 170, C(0)                                                                                                                                                                                                                                                                                                                                                                   |
| 230 | 900 | W230 DATA | @_UINT/CC/SCALbx34_ARA0 te=230-te-230 write args=0, 25, Cu(1859660671);@_SINT/CC/SCALbx16_ARA0 te=230-te-230 write args=0, 169, C(-3)                                                                                                                                                                                                                                                                                                                                                                  |
| 231 | 900 | W231 DATA | @_UINT/CC/SCALbx34_ARA0 te=231-te-231 write args=0, 24, Cu(1780037320);@_SINT/CC/SCALbx16_ARA0 te=231-te-231 write args=0, 168, C(5)                                                                                                                                                                                                                                                                                                                                                                   |
| 232 | 900 | W232 DATA | @_UINT/CC/SCALbx34_ARA0 te=232-te-232 write args=0, 23, Cu(1381403509);@_SINT/CC/SCALbx16_ARA0 te=232-te-232 write args=0, 167, C(-2)                                                                                                                                                                                                                                                                                                                                                                  |
| 233 | 900 | W233 DATA | @_UINT/CC/SCALbx34_ARA0 te=233-te-233 write args=0, 22, Cu(1452775106);@_SINT/CC/SCALbx16_ARA0 te=233-te-233 write args=0, 166, C(0)                                                                                                                                                                                                                                                                                                                                                                   |
| 234 | 900 | W234 DATA | @_UINT/CC/SCALbx34_ARA0 te=234-te-234 write args=0, 21, Cu(1540665371);@_SINT/CC/SCALbx16_ARA0 te=234-te-234 write args=0, 165, C(-2)                                                                                                                                                                                                                                                                                                                                                                  |
| 235 | 900 | W235 DATA | @_UINT/CC/SCALbx34_ARA0 te=235-te-235 write args=0, 20, Cu(1595256236);@_SINT/CC/SCALbx16_ARA0 te=235-te-235 write args=0, 164, C(-5)                                                                                                                                                                                                                                                                                                                                                                  |
| 236 | 900 | W236 DATA | @_UINT/CC/SCALbx34_ARA0 te=236-te-236 write args=0, 19, Cu(1095957929);@_SINT/CC/SCALbx16_ARA0 te=236-te-236 write args=0, 163, C(0)                                                                                                                                                                                                                                                                                                                                                                   |
| 237 | 900 | W237 DATA | @_UINT/CC/SCALbx34_ARA0 te=237-te-237 write args=0, 18, Cu(1167319070);@_SINT/CC/SCALbx16_ARA0 te=237-te-237 write args=0, 162, C(0)                                                                                                                                                                                                                                                                                                                                                                   |
| 238 | 900 | W238 DATA | @_UINT/CC/SCALbx34_ARA0 te=238-te-238 write args=0, 17, Cu(1221641927);@_SINT/CC/SCALbx16_ARA0 te=238-te-238 write args=0, 161, C(-5)                                                                                                                                                                                                                                                                                                                                                                  |
| 239 | 900 | W239 DATA | @_UINT/CC/SCALbx34_ARA0 te=239-te-239 write args=0, 16, Cu(1276238704);@_SINT/CC/SCALbx16_ARA0 te=239-te-239 write args=0, 160, C(-1)                                                                                                                                                                                                                                                                                                                                                                  |
| 240 | 900 | W240 DATA | @_UINT/CC/SCALbx34_ARA0 te=240-te-240 write args=0, 15, Cu(944750013);@_SINT/CC/SCALbx16_ARA0 te=240-te-240 write args=0, 159, C(-1)                                                                                                                                                                                                                                                                                                                                                                   |
| 241 | 900 | W241 DATA | @_UINT/CC/SCALbx34_ARA0 te=241-te-241 write args=0, 14, Cu(1015980042);@_SINT/CC/SCALbx16_ARA0 te=241-te-241 write args=0, 158, C(-5)                                                                                                                                                                                                                                                                                                                                                                  |
| 242 | 900 | W242 DATA | @_UINT/CC/SCALbx34_ARA0 te=242-te-242 write args=0, 13, Cu(835552979);@_SINT/CC/SCALbx16_ARA0 te=242-te-242 write args=0, 157, C(4)                                                                                                                                                                                                                                                                                                                                                                    |
| 243 | 900 | W243 DATA | @_UINT/CC/SCALbx34_ARA0 te=243-te-243 write args=0, 12, Cu(890018660);@_SINT/CC/SCALbx16_ARA0 te=243-te-243 write args=0, 156, C(0)                                                                                                                                                                                                                                                                                                                                                                    |
| 244 | 900 | W244 DATA | @_UINT/CC/SCALbx34_ARA0 te=244-te-244 write args=0, 11, Cu(726387553);@_SINT/CC/SCALbx16_ARA0 te=244-te-244 write args=0, 155, C(-1)                                                                                                                                                                                                                                                                                                                                                                   |
| 245 | 900 | W245 DATA | @_UINT/CC/SCALbx34_ARA0 te=245-te-245 write args=0, 10, Cu(797628118);@_SINT/CC/SCALbx16_ARA0 te=245-te-245 write args=0, 154, C(-2)                                                                                                                                                                                                                                                                                                                                                                   |
| 246 | 900 | W246 DATA | @_UINT/CC/SCALbx34_ARA0 te=246-te-246 write args=0, 9, Cu(583659535);@_SINT/CC/SCALbx16_ARA0 te=246-te-246 write args=0, 153, C(-2)                                                                                                                                                                                                                                                                                                                                                                    |
| 247 | 900 | W247 DATA | @_UINT/CC/SCALbx34_ARA0 te=247-te-247 write args=0, 8, Cu(638119352);@_SINT/CC/SCALbx16_ARA0 te=247-te-247 write args=0, 152, C(-2)                                                                                                                                                                                                                                                                                                                                                                    |
| 248 | 900 | W248 DATA | @_UINT/CC/SCALbx34_ARA0 te=248-te-248 write args=0, 7, Cu(507990021);@_SINT/CC/SCALbx16_ARA0 te=248-te-248 write args=0, 151, C(-2)                                                                                                                                                                                                                                                                                                                                                                    |
| 249 | 900 | W249 DATA | @_UINT/CC/SCALbx34_ARA0 te=249-te-249 write args=0, 6, Cu(445009330);@_SINT/CC/SCALbx16_ARA0 te=249-te-249 write args=0, 150, C(2)                                                                                                                                                                                                                                                                                                                                                                     |
| 250 | 900 | W250 DATA | @_UINT/CC/SCALbx34_ARA0 te=250-te-250 write args=0, 5, Cu(398814059);@_SINT/CC/SCALbx16_ARA0 te=250-te-250 write args=0, 149, C(2)                                                                                                                                                                                                                                                                                                                                                                     |
| 251 | 900 | W251 DATA | @_UINT/CC/SCALbx34_ARA0 te=251-te-251 write args=0, 4, Cu(319059676);@_SINT/CC/SCALbx16_ARA0 te=251-te-251 write args=0, 148, C(-2)                                                                                                                                                                                                                                                                                                                                                                    |
| 252 | 900 | W252 DATA | @_UINT/CC/SCALbx34_ARA0 te=252-te-252 write args=0, 3, Cu(222504665);@_SINT/CC/SCALbx16_ARA0 te=252-te-252 write args=0, 147, C(5)                                                                                                                                                                                                                                                                                                                                                                     |
| 253 | 900 | W253 DATA | @_UINT/CC/SCALbx34_ARA0 te=253-te-253 write args=0, 2, Cu(159529838);@_SINT/CC/SCALbx16_ARA0 te=253-te-253 write args=0, 146, C(-2)                                                                                                                                                                                                                                                                                                                                                                    |
| 254 | 900 | W254 DATA | @_UINT/CC/SCALbx34_ARA0 te=254-te-254 write args=0, 1, Cu(79764919);@_SINT/CC/SCALbx16_ARA0 te=254-te-254 write args=0, 145, C(-3)                                                                                                                                                                                                                                                                                                                                                                     |
| 255 | 900 | W255 DATA | @_UINT/CC/SCALbx34_ARA0 te=255-te-255 write args=0, 0, Cu(0);@_SINT/CC/SCALbx16_ARA0 te=255-te-255 write args=0, 144, C(1)                                                                                                                                                                                                                                                                                                                                                                             |
| 256 | 900 | W256 DATA | @_SINT/CC/SCALbx16_ARA0 te=256-te-256 write args=0, 143, C(-2)                                                                                                                                                                                                                                                                                                                                                                                                                                         |
| 257 | 900 | W257 DATA | @_SINT/CC/SCALbx16_ARA0 te=257-te-257 write args=0, 142, C(-2)                                                                                                                                                                                                                                                                                                                                                                                                                                         |
| 258 | 900 | W258 DATA | @_SINT/CC/SCALbx16_ARA0 te=258-te-258 write args=0, 141, C(-2)                                                                                                                                                                                                                                                                                                                                                                                                                                         |
| 259 | 900 | W259 DATA | @_SINT/CC/SCALbx16_ARA0 te=259-te-259 write args=0, 140, C(-1)                                                                                                                                                                                                                                                                                                                                                                                                                                         |
| 260 | 900 | W260 DATA | @_SINT/CC/SCALbx16_ARA0 te=260-te-260 write args=0, 139, C(0)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 261 | 900 | W261 DATA | @_SINT/CC/SCALbx16_ARA0 te=261-te-261 write args=0, 138, C(-3)                                                                                                                                                                                                                                                                                                                                                                                                                                         |
| 262 | 900 | W262 DATA | @_SINT/CC/SCALbx16_ARA0 te=262-te-262 write args=0, 137, C(-2)                                                                                                                                                                                                                                                                                                                                                                                                                                         |
| 263 | 900 | W263 DATA | @_SINT/CC/SCALbx16_ARA0 te=263-te-263 write args=0, 136, C(-1)                                                                                                                                                                                                                                                                                                                                                                                                                                         |
| 264 | 900 | W264 DATA | @_SINT/CC/SCALbx16_ARA0 te=264-te-264 write args=0, 135, C(-1)                                                                                                                                                                                                                                                                                                                                                                                                                                         |
| 265 | 900 | W265 DATA | @_SINT/CC/SCALbx16_ARA0 te=265-te-265 write args=0, 134, C(2)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 266 | 900 | W266 DATA | @_SINT/CC/SCALbx16_ARA0 te=266-te-266 write args=0, 133, C(3)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 267 | 900 | W267 DATA | @_SINT/CC/SCALbx16_ARA0 te=267-te-267 write args=0, 132, C(0)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 268 | 900 | W268 DATA | @_SINT/CC/SCALbx16_ARA0 te=268-te-268 write args=0, 131, C(2)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 269 | 900 | W269 DATA | @_SINT/CC/SCALbx16_ARA0 te=269-te-269 write args=0, 130, C(-2)                                                                                                                                                                                                                                                                                                                                                                                                                                         |
| 270 | 900 | W270 DATA | @_SINT/CC/SCALbx16_ARA0 te=270-te-270 write args=0, 129, C(-2)                                                                                                                                                                                                                                                                                                                                                                                                                                         |
| 271 | 900 | W271 DATA | @_SINT/CC/SCALbx16_ARA0 te=271-te-271 write args=0, 128, C(0)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 272 | 900 | W272 DATA | @_SINT/CC/SCALbx16_ARA0 te=272-te-272 write args=0, 127, C(-2)                                                                                                                                                                                                                                                                                                                                                                                                                                         |
| 273 | 900 | W273 DATA | @_SINT/CC/SCALbx16_ARA0 te=273-te-273 write args=0, 126, C(6)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 274 | 900 | W274 DATA | @_SINT/CC/SCALbx16_ARA0 te=274-te-274 write args=0, 125, C(-2)                                                                                                                                                                                                                                                                                                                                                                                                                                         |
| 275 | 900 | W275 DATA | @_SINT/CC/SCALbx16_ARA0 te=275-te-275 write args=0, 124, C(-2)                                                                                                                                                                                                                                                                                                                                                                                                                                         |
| 276 | 900 | W276 DATA | @_SINT/CC/SCALbx16_ARA0 te=276-te-276 write args=0, 123, C(1)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 277 | 900 | W277 DATA | @_SINT/CC/SCALbx16_ARA0 te=277-te-277 write args=0, 122, C(1)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 278 | 900 | W278 DATA | @_SINT/CC/SCALbx16_ARA0 te=278-te-278 write args=0, 121, C(-3)                                                                                                                                                                                                                                                                                                                                                                                                                                         |
| 279 | 900 | W279 DATA | @_SINT/CC/SCALbx16_ARA0 te=279-te-279 write args=0, 120, C(-1)                                                                                                                                                                                                                                                                                                                                                                                                                                         |
| 280 | 900 | W280 DATA | @_SINT/CC/SCALbx16_ARA0 te=280-te-280 write args=0, 119, C(-5)                                                                                                                                                                                                                                                                                                                                                                                                                                         |
| 281 | 900 | W281 DATA | @_SINT/CC/SCALbx16_ARA0 te=281-te-281 write args=0, 118, C(-7)                                                                                                                                                                                                                                                                                                                                                                                                                                         |
| 282 | 900 | W282 DATA | @_SINT/CC/SCALbx16_ARA0 te=282-te-282 write args=0, 117, C(-1)                                                                                                                                                                                                                                                                                                                                                                                                                                         |
| 283 | 900 | W283 DATA | @_SINT/CC/SCALbx16_ARA0 te=283-te-283 write args=0, 116, C(0)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 284 | 900 | W284 DATA | @_SINT/CC/SCALbx16_ARA0 te=284-te-284 write args=0, 115, C(1)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 285 | 900 | W285 DATA | @_SINT/CC/SCALbx16_ARA0 te=285-te-285 write args=0, 114, C(-3)                                                                                                                                                                                                                                                                                                                                                                                                                                         |
| 286 | 900 | W286 DATA | @_SINT/CC/SCALbx16_ARA0 te=286-te-286 write args=0, 113, C(-1)                                                                                                                                                                                                                                                                                                                                                                                                                                         |
| 287 | 900 | W287 DATA | @_SINT/CC/SCALbx16_ARA0 te=287-te-287 write args=0, 112, C(-1)                                                                                                                                                                                                                                                                                                                                                                                                                                         |
| 288 | 900 | W288 DATA | @_SINT/CC/SCALbx16_ARA0 te=288-te-288 write args=0, 111, C(0)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 289 | 900 | W289 DATA | @_SINT/CC/SCALbx16_ARA0 te=289-te-289 write args=0, 110, C(-3)                                                                                                                                                                                                                                                                                                                                                                                                                                         |
| 290 | 900 | W290 DATA | @_SINT/CC/SCALbx16_ARA0 te=290-te-290 write args=0, 109, C(-4)                                                                                                                                                                                                                                                                                                                                                                                                                                         |
| 291 | 900 | W291 DATA | @_SINT/CC/SCALbx16_ARA0 te=291-te-291 write args=0, 108, C(-2)                                                                                                                                                                                                                                                                                                                                                                                                                                         |
| 292 | 900 | W292 DATA | @_SINT/CC/SCALbx16_ARA0 te=292-te-292 write args=0, 107, C(-3)                                                                                                                                                                                                                                                                                                                                                                                                                                         |
| 293 | 900 | W293 DATA | @_SINT/CC/SCALbx16_ARA0 te=293-te-293 write args=0, 106, C(-2)                                                                                                                                                                                                                                                                                                                                                                                                                                         |
| 294 | 900 | W294 DATA | @_SINT/CC/SCALbx16_ARA0 te=294-te-294 write args=0, 105, C(5)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 295 | 900 | W295 DATA | @_SINT/CC/SCALbx16_ARA0 te=295-te-295 write args=0, 104, C(-5)                                                                                                                                                                                                                                                                                                                                                                                                                                         |
| 296 | 900 | W296 DATA | @_SINT/CC/SCALbx16_ARA0 te=296-te-296 write args=0, 103, C(0)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 297 | 900 | W297 DATA | @_SINT/CC/SCALbx16_ARA0 te=297-te-297 write args=0, 102, C(1)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 298 | 900 | W298 DATA | @_SINT/CC/SCALbx16_ARA0 te=298-te-298 write args=0, 101, C(-3)                                                                                                                                                                                                                                                                                                                                                                                                                                         |
| 299 | 900 | W299 DATA | @_SINT/CC/SCALbx16_ARA0 te=299-te-299 write args=0, 100, C(1)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 300 | 900 | W300 DATA | @_SINT/CC/SCALbx16_ARA0 te=300-te-300 write args=0, 99, C(7)                                                                                                                                                                                                                                                                                                                                                                                                                                           |
| 301 | 900 | W301 DATA | @_SINT/CC/SCALbx16_ARA0 te=301-te-301 write args=0, 98, C(0)                                                                                                                                                                                                                                                                                                                                                                                                                                           |
| 302 | 900 | W302 DATA | @_SINT/CC/SCALbx16_ARA0 te=302-te-302 write args=0, 97, C(-1)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 303 | 900 | W303 DATA | @_SINT/CC/SCALbx16_ARA0 te=303-te-303 write args=0, 96, C(-3)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 304 | 900 | W304 DATA | @_SINT/CC/SCALbx16_ARA0 te=304-te-304 write args=0, 95, C(-3)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 305 | 900 | W305 DATA | @_SINT/CC/SCALbx16_ARA0 te=305-te-305 write args=0, 94, C(-4)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 306 | 900 | W306 DATA | @_SINT/CC/SCALbx16_ARA0 te=306-te-306 write args=0, 93, C(-5)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 307 | 900 | W307 DATA | @_SINT/CC/SCALbx16_ARA0 te=307-te-307 write args=0, 92, C(-5)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 308 | 900 | W308 DATA | @_SINT/CC/SCALbx16_ARA0 te=308-te-308 write args=0, 91, C(-4)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 309 | 900 | W309 DATA | @_SINT/CC/SCALbx16_ARA0 te=309-te-309 write args=0, 90, C(0)                                                                                                                                                                                                                                                                                                                                                                                                                                           |
| 310 | 900 | W310 DATA | @_SINT/CC/SCALbx16_ARA0 te=310-te-310 write args=0, 89, C(2)                                                                                                                                                                                                                                                                                                                                                                                                                                           |
| 311 | 900 | W311 DATA | @_SINT/CC/SCALbx16_ARA0 te=311-te-311 write args=0, 88, C(-5)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 312 | 900 | W312 DATA | @_SINT/CC/SCALbx16_ARA0 te=312-te-312 write args=0, 87, C(1)                                                                                                                                                                                                                                                                                                                                                                                                                                           |
| 313 | 900 | W313 DATA | @_SINT/CC/SCALbx16_ARA0 te=313-te-313 write args=0, 86, C(-2)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 314 | 900 | W314 DATA | @_SINT/CC/SCALbx16_ARA0 te=314-te-314 write args=0, 85, C(-5)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 315 | 900 | W315 DATA | @_SINT/CC/SCALbx16_ARA0 te=315-te-315 write args=0, 84, C(9)                                                                                                                                                                                                                                                                                                                                                                                                                                           |
| 316 | 900 | W316 DATA | @_SINT/CC/SCALbx16_ARA0 te=316-te-316 write args=0, 83, C(-5)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 317 | 900 | W317 DATA | @_SINT/CC/SCALbx16_ARA0 te=317-te-317 write args=0, 82, C(-6)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 318 | 900 | W318 DATA | @_SINT/CC/SCALbx16_ARA0 te=318-te-318 write args=0, 81, C(-4)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 319 | 900 | W319 DATA | @_SINT/CC/SCALbx16_ARA0 te=319-te-319 write args=0, 80, C(-4)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 320 | 900 | W320 DATA | @_SINT/CC/SCALbx16_ARA0 te=320-te-320 write args=0, 79, C(-4)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 321 | 900 | W321 DATA | @_SINT/CC/SCALbx16_ARA0 te=321-te-321 write args=0, 78, C(-7)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 322 | 900 | W322 DATA | @_SINT/CC/SCALbx16_ARA0 te=322-te-322 write args=0, 77, C(-2)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 323 | 900 | W323 DATA | @_SINT/CC/SCALbx16_ARA0 te=323-te-323 write args=0, 76, C(0)                                                                                                                                                                                                                                                                                                                                                                                                                                           |
| 324 | 900 | W324 DATA | @_SINT/CC/SCALbx16_ARA0 te=324-te-324 write args=0, 75, C(0)                                                                                                                                                                                                                                                                                                                                                                                                                                           |
| 325 | 900 | W325 DATA | @_SINT/CC/SCALbx16_ARA0 te=325-te-325 write args=0, 74, C(-1)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 326 | 900 | W326 DATA | @_SINT/CC/SCALbx16_ARA0 te=326-te-326 write args=0, 73, C(2)                                                                                                                                                                                                                                                                                                                                                                                                                                           |
| 327 | 900 | W327 DATA | @_SINT/CC/SCALbx16_ARA0 te=327-te-327 write args=0, 72, C(-1)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 328 | 900 | W328 DATA | @_SINT/CC/SCALbx16_ARA0 te=328-te-328 write args=0, 71, C(1)                                                                                                                                                                                                                                                                                                                                                                                                                                           |
| 329 | 900 | W329 DATA | @_SINT/CC/SCALbx16_ARA0 te=329-te-329 write args=0, 70, C(-2)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 330 | 900 | W330 DATA | @_SINT/CC/SCALbx16_ARA0 te=330-te-330 write args=0, 69, C(-3)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 331 | 900 | W331 DATA | @_SINT/CC/SCALbx16_ARA0 te=331-te-331 write args=0, 68, C(0)                                                                                                                                                                                                                                                                                                                                                                                                                                           |
| 332 | 900 | W332 DATA | @_SINT/CC/SCALbx16_ARA0 te=332-te-332 write args=0, 67, C(-2)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 333 | 900 | W333 DATA | @_SINT/CC/SCALbx16_ARA0 te=333-te-333 write args=0, 66, C(1)                                                                                                                                                                                                                                                                                                                                                                                                                                           |
| 334 | 900 | W334 DATA | @_SINT/CC/SCALbx16_ARA0 te=334-te-334 write args=0, 65, C(0)                                                                                                                                                                                                                                                                                                                                                                                                                                           |
| 335 | 900 | W335 DATA | @_SINT/CC/SCALbx16_ARA0 te=335-te-335 write args=0, 64, C(-5)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 336 | 900 | W336 DATA | @_SINT/CC/SCALbx16_ARA0 te=336-te-336 write args=0, 63, C(4)                                                                                                                                                                                                                                                                                                                                                                                                                                           |
| 337 | 900 | W337 DATA | @_SINT/CC/SCALbx16_ARA0 te=337-te-337 write args=0, 62, C(3)                                                                                                                                                                                                                                                                                                                                                                                                                                           |
| 338 | 900 | W338 DATA | @_SINT/CC/SCALbx16_ARA0 te=338-te-338 write args=0, 61, C(-5)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 339 | 900 | W339 DATA | @_SINT/CC/SCALbx16_ARA0 te=339-te-339 write args=0, 60, C(0)                                                                                                                                                                                                                                                                                                                                                                                                                                           |
| 340 | 900 | W340 DATA | @_SINT/CC/SCALbx16_ARA0 te=340-te-340 write args=0, 59, C(-4)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 341 | 900 | W341 DATA | @_SINT/CC/SCALbx16_ARA0 te=341-te-341 write args=0, 58, C(-7)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 342 | 900 | W342 DATA | @_SINT/CC/SCALbx16_ARA0 te=342-te-342 write args=0, 57, C(-2)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 343 | 900 | W343 DATA | @_SINT/CC/SCALbx16_ARA0 te=343-te-343 write args=0, 56, C(0)                                                                                                                                                                                                                                                                                                                                                                                                                                           |
| 344 | 900 | W344 DATA | @_SINT/CC/SCALbx16_ARA0 te=344-te-344 write args=0, 55, C(0)                                                                                                                                                                                                                                                                                                                                                                                                                                           |
| 345 | 900 | W345 DATA | @_SINT/CC/SCALbx16_ARA0 te=345-te-345 write args=0, 54, C(-1)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 346 | 900 | W346 DATA | @_SINT/CC/SCALbx16_ARA0 te=346-te-346 write args=0, 53, C(2)                                                                                                                                                                                                                                                                                                                                                                                                                                           |
| 347 | 900 | W347 DATA | @_SINT/CC/SCALbx16_ARA0 te=347-te-347 write args=0, 52, C(-1)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 348 | 900 | W348 DATA | @_SINT/CC/SCALbx16_ARA0 te=348-te-348 write args=0, 51, C(2)                                                                                                                                                                                                                                                                                                                                                                                                                                           |
| 349 | 900 | W349 DATA | @_SINT/CC/SCALbx16_ARA0 te=349-te-349 write args=0, 50, C(-3)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 350 | 900 | W350 DATA | @_SINT/CC/SCALbx16_ARA0 te=350-te-350 write args=0, 49, C(-4)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 351 | 900 | W351 DATA | @_SINT/CC/SCALbx16_ARA0 te=351-te-351 write args=0, 48, C(0)                                                                                                                                                                                                                                                                                                                                                                                                                                           |
| 352 | 900 | W352 DATA | @_SINT/CC/SCALbx16_ARA0 te=352-te-352 write args=0, 47, C(-2)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 353 | 900 | W353 DATA | @_SINT/CC/SCALbx16_ARA0 te=353-te-353 write args=0, 46, C(1)                                                                                                                                                                                                                                                                                                                                                                                                                                           |
| 354 | 900 | W354 DATA | @_SINT/CC/SCALbx16_ARA0 te=354-te-354 write args=0, 45, C(1)                                                                                                                                                                                                                                                                                                                                                                                                                                           |
| 355 | 900 | W355 DATA | @_SINT/CC/SCALbx16_ARA0 te=355-te-355 write args=0, 44, C(-6)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 356 | 900 | W356 DATA | @_SINT/CC/SCALbx16_ARA0 te=356-te-356 write args=0, 43, C(3)                                                                                                                                                                                                                                                                                                                                                                                                                                           |
| 357 | 900 | W357 DATA | @_SINT/CC/SCALbx16_ARA0 te=357-te-357 write args=0, 42, C(4)                                                                                                                                                                                                                                                                                                                                                                                                                                           |
| 358 | 900 | W358 DATA | @_SINT/CC/SCALbx16_ARA0 te=358-te-358 write args=0, 41, C(-5)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 359 | 900 | W359 DATA | @_SINT/CC/SCALbx16_ARA0 te=359-te-359 write args=0, 40, C(0)                                                                                                                                                                                                                                                                                                                                                                                                                                           |
| 360 | 900 | W360 DATA | @_SINT/CC/SCALbx16_ARA0 te=360-te-360 write args=0, 39, C(0)                                                                                                                                                                                                                                                                                                                                                                                                                                           |
| 361 | 900 | W361 DATA | @_SINT/CC/SCALbx16_ARA0 te=361-te-361 write args=0, 38, C(-8)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 362 | 900 | W362 DATA | @_SINT/CC/SCALbx16_ARA0 te=362-te-362 write args=0, 37, C(-2)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 363 | 900 | W363 DATA | @_SINT/CC/SCALbx16_ARA0 te=363-te-363 write args=0, 36, C(-2)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 364 | 900 | W364 DATA | @_SINT/CC/SCALbx16_ARA0 te=364-te-364 write args=0, 35, C(0)                                                                                                                                                                                                                                                                                                                                                                                                                                           |
| 365 | 900 | W365 DATA | @_SINT/CC/SCALbx16_ARA0 te=365-te-365 write args=0, 34, C(-4)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 366 | 900 | W366 DATA | @_SINT/CC/SCALbx16_ARA0 te=366-te-366 write args=0, 33, C(-5)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 367 | 900 | W367 DATA | @_SINT/CC/SCALbx16_ARA0 te=367-te-367 write args=0, 32, C(-3)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 368 | 900 | W368 DATA | @_SINT/CC/SCALbx16_ARA0 te=368-te-368 write args=0, 31, C(-4)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 369 | 900 | W369 DATA | @_SINT/CC/SCALbx16_ARA0 te=369-te-369 write args=0, 30, C(-5)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 370 | 900 | W370 DATA | @_SINT/CC/SCALbx16_ARA0 te=370-te-370 write args=0, 29, C(-6)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 371 | 900 | W371 DATA | @_SINT/CC/SCALbx16_ARA0 te=371-te-371 write args=0, 28, C(-5)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 372 | 900 | W372 DATA | @_SINT/CC/SCALbx16_ARA0 te=372-te-372 write args=0, 27, C(-2)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 373 | 900 | W373 DATA | @_SINT/CC/SCALbx16_ARA0 te=373-te-373 write args=0, 26, C(-3)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 374 | 900 | W374 DATA | @_SINT/CC/SCALbx16_ARA0 te=374-te-374 write args=0, 25, C(-3)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 375 | 900 | W375 DATA | @_SINT/CC/SCALbx16_ARA0 te=375-te-375 write args=0, 24, C(-4)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 376 | 900 | W376 DATA | @_SINT/CC/SCALbx16_ARA0 te=376-te-376 write args=0, 23, C(-5)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 377 | 900 | W377 DATA | @_SINT/CC/SCALbx16_ARA0 te=377-te-377 write args=0, 22, C(-5)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 378 | 900 | W378 DATA | @_SINT/CC/SCALbx16_ARA0 te=378-te-378 write args=0, 21, C(12)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 379 | 900 | W379 DATA | @_SINT/CC/SCALbx16_ARA0 te=379-te-379 write args=0, 20, C(-2)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 380 | 900 | W380 DATA | @_SINT/CC/SCALbx16_ARA0 te=380-te-380 write args=0, 19, C(-3)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 381 | 900 | W381 DATA | @_SINT/CC/SCALbx16_ARA0 te=381-te-381 write args=0, 18, C(-1)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 382 | 900 | W382 DATA | @_SINT/CC/SCALbx16_ARA0 te=382-te-382 write args=0, 17, C(0)                                                                                                                                                                                                                                                                                                                                                                                                                                           |
| 383 | 900 | W383 DATA | @_SINT/CC/SCALbx16_ARA0 te=383-te-383 write args=0, 16, C(1)                                                                                                                                                                                                                                                                                                                                                                                                                                           |
| 384 | 900 | W384 DATA | @_SINT/CC/SCALbx16_ARA0 te=384-te-384 write args=0, 15, C(1)                                                                                                                                                                                                                                                                                                                                                                                                                                           |
| 385 | 900 | W385 DATA | @_SINT/CC/SCALbx16_ARA0 te=385-te-385 write args=0, 14, C(-2)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 386 | 900 | W386 DATA | @_SINT/CC/SCALbx16_ARA0 te=386-te-386 write args=0, 13, C(0)                                                                                                                                                                                                                                                                                                                                                                                                                                           |
| 387 | 900 | W387 DATA | @_SINT/CC/SCALbx16_ARA0 te=387-te-387 write args=0, 12, C(1)                                                                                                                                                                                                                                                                                                                                                                                                                                           |
| 388 | 900 | W388 DATA | @_SINT/CC/SCALbx16_ARA0 te=388-te-388 write args=0, 11, C(0)                                                                                                                                                                                                                                                                                                                                                                                                                                           |
| 389 | 900 | W389 DATA | @_SINT/CC/SCALbx16_ARA0 te=389-te-389 write args=0, 10, C(-1)                                                                                                                                                                                                                                                                                                                                                                                                                                          |
| 390 | 900 | W390 DATA | @_SINT/CC/SCALbx16_ARA0 te=390-te-390 write args=0, 9, C(-2)                                                                                                                                                                                                                                                                                                                                                                                                                                           |
| 391 | 900 | W391 DATA | @_SINT/CC/SCALbx16_ARA0 te=391-te-391 write args=0, 8, C(-1)                                                                                                                                                                                                                                                                                                                                                                                                                                           |
| 392 | 900 | W392 DATA | @_SINT/CC/SCALbx16_ARA0 te=392-te-392 write args=0, 7, C(-1)                                                                                                                                                                                                                                                                                                                                                                                                                                           |
| 393 | 900 | W393 DATA | @_SINT/CC/SCALbx16_ARA0 te=393-te-393 write args=0, 6, C(-1)                                                                                                                                                                                                                                                                                                                                                                                                                                           |
| 394 | 900 | W394 DATA | @_SINT/CC/SCALbx16_ARA0 te=394-te-394 write args=0, 5, C(1)                                                                                                                                                                                                                                                                                                                                                                                                                                            |
| 395 | 900 | W395 DATA | @_SINT/CC/SCALbx16_ARA0 te=395-te-395 write args=0, 4, C(-4)                                                                                                                                                                                                                                                                                                                                                                                                                                           |
| 396 | 900 | W396 DATA | @_SINT/CC/SCALbx16_ARA0 te=396-te-396 write args=0, 3, C(0)                                                                                                                                                                                                                                                                                                                                                                                                                                            |
| 397 | 900 | W397 DATA | @_SINT/CC/SCALbx16_ARA0 te=397-te-397 write args=0, 2, C(0)                                                                                                                                                                                                                                                                                                                                                                                                                                            |
| 398 | 900 | W398 DATA | @_SINT/CC/SCALbx16_ARA0 te=398-te-398 write args=0, 1, C(-2)                                                                                                                                                                                                                                                                                                                                                                                                                                           |
| 399 | 900 | W399 DATA | @_SINT/CC/SCALbx16_ARA0 te=399-te-399 write args=0, 0, C(2)                                                                                                                                                                                                                                                                                                                                                                                                                                            |
| 400 | 900 | W400 DATA |                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        |
*-----+-----+-----------+--------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------*

// Restructure Technology Settings
*------------------------+---------+---------------------------------------------------------------------------------*
| Key                    | Value   | Description                                                                     |
*------------------------+---------+---------------------------------------------------------------------------------*
| int_flr_mul            | 16000   |                                                                                 |
| fp_fl_dp_div           | 5       |                                                                                 |
| fp_fl_dp_add           | 5       |                                                                                 |
| fp_fl_dp_mul           | 5       |                                                                                 |
| fp_fl_sp_div           | 5       |                                                                                 |
| fp_fl_sp_add           | 5       |                                                                                 |
| fp_fl_sp_mul           | 5       |                                                                                 |
| max_no_fp_muls         | 6       | Maximum number of adders and subtractors (or combos) to instantiate per thread. |
| max_no_fp_muls         | 6       | Maximum number of f/p dividers to instantiate per thread.                       |
| max_no_int_muls        | 3       | Maximum number of int multipliers to instantiate per thread.                    |
| max_no_fp_divs         | 2       | Maximum number of f/p dividers to instantiate per thread.                       |
| max_no_int_divs        | 2       | Maximum number of int dividers to instantiate per thread.                       |
| res2-offchip-threshold | 1000000 |                                                                                 |
| res2-combram-threshold | 32      |                                                                                 |
| res2-regfile-threshold | 8       |                                                                                 |
*------------------------+---------+---------------------------------------------------------------------------------*

// Offchip Memory Physical Ports/Banks
*-----------+----------+----------+--------+--------+-------+-----------*
| Name      | Protocol | No Words | Awidth | Dwidth | Lanes | LaneWidth |
*-----------+----------+----------+--------+--------+-------+-----------*
| dram0bank | HFAST1   | 4194304  | 22     | 256    | 32    | 8         |
*-----------+----------+----------+--------+--------+-------+-----------*

// */

//  
// LCP delay estimations included: turn off with -vnl-lcp-delay-estimate=disable
// eof (HPR L/S Verilog)
